magic
tech sky130A
magscale 1 2
timestamp 1700843682
<< obsli1 >>
rect 1104 2159 9016 9809
<< obsm1 >>
rect 14 1708 9094 9840
<< metal2 >>
rect 5814 11556 5870 12356
rect 18 0 74 800
rect 8390 0 8446 800
<< obsm2 >>
rect 20 11500 5758 11556
rect 5926 11500 9090 11556
rect 20 856 9090 11500
rect 130 800 8334 856
rect 8502 800 9090 856
<< metal3 >>
rect 0 8848 800 8968
rect 9412 7488 10212 7608
<< obsm3 >>
rect 800 9048 9412 9825
rect 880 8768 9412 9048
rect 800 7688 9412 8768
rect 800 7408 9332 7688
rect 800 2143 9412 7408
<< metal4 >>
rect 1933 2128 2253 9840
rect 2593 2128 2913 9840
rect 3911 2128 4231 9840
rect 4571 2128 4891 9840
rect 5889 2128 6209 9840
rect 6549 2128 6869 9840
rect 7867 2128 8187 9840
rect 8527 2128 8847 9840
<< metal5 >>
rect 1056 9340 9064 9660
rect 1056 8680 9064 9000
rect 1056 7436 9064 7756
rect 1056 6776 9064 7096
rect 1056 5532 9064 5852
rect 1056 4872 9064 5192
rect 1056 3628 9064 3948
rect 1056 2968 9064 3288
<< labels >>
rlabel metal4 s 2593 2128 2913 9840 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 4571 2128 4891 9840 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 6549 2128 6869 9840 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 8527 2128 8847 9840 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 3628 9064 3948 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 5532 9064 5852 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 7436 9064 7756 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 9340 9064 9660 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 1933 2128 2253 9840 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 3911 2128 4231 9840 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 5889 2128 6209 9840 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 7867 2128 8187 9840 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 2968 9064 3288 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 4872 9064 5192 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 6776 9064 7096 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 8680 9064 9000 6 VPWR
port 2 nsew power bidirectional
rlabel metal3 s 0 8848 800 8968 6 clk
port 3 nsew signal input
rlabel metal2 s 18 0 74 800 6 clkout
port 4 nsew signal output
rlabel metal3 s 9412 7488 10212 7608 6 reset
port 5 nsew signal input
rlabel metal2 s 5814 11556 5870 12356 6 sel[0]
port 6 nsew signal input
rlabel metal2 s 8390 0 8446 800 6 sel[1]
port 7 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 10212 12356
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 822622
string GDS_FILE /home/rohith_nagesh/Baud-rate-generator/openlane/pes_brg/runs/23_11_24_22_02/results/signoff/pes_brg.magic.gds
string GDS_START 429172
<< end >>

