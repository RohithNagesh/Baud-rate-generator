magic
tech sky130A
magscale 1 2
timestamp 1700843680
<< viali >>
rect 2421 9673 2455 9707
rect 5549 9673 5583 9707
rect 5917 9673 5951 9707
rect 3433 9605 3467 9639
rect 1593 9537 1627 9571
rect 3341 9537 3375 9571
rect 3617 9537 3651 9571
rect 4077 9517 4111 9551
rect 4537 9537 4571 9571
rect 5733 9537 5767 9571
rect 6101 9537 6135 9571
rect 6469 9537 6503 9571
rect 6561 9537 6595 9571
rect 6837 9537 6871 9571
rect 7564 9537 7598 9571
rect 1961 9469 1995 9503
rect 2053 9469 2087 9503
rect 2145 9469 2179 9503
rect 2237 9469 2271 9503
rect 2513 9469 2547 9503
rect 3985 9469 4019 9503
rect 4353 9469 4387 9503
rect 4445 9469 4479 9503
rect 6745 9469 6779 9503
rect 7297 9469 7331 9503
rect 3157 9401 3191 9435
rect 3617 9401 3651 9435
rect 1777 9333 1811 9367
rect 3801 9333 3835 9367
rect 4721 9333 4755 9367
rect 7021 9333 7055 9367
rect 8677 9333 8711 9367
rect 5825 9129 5859 9163
rect 4261 9061 4295 9095
rect 2881 8993 2915 9027
rect 5641 8993 5675 9027
rect 3157 8925 3191 8959
rect 3249 8925 3283 8959
rect 3479 8925 3513 8959
rect 3617 8925 3651 8959
rect 7113 8925 7147 8959
rect 7389 8925 7423 8959
rect 7665 8925 7699 8959
rect 7849 8925 7883 8959
rect 8401 8925 8435 8959
rect 8493 8925 8527 8959
rect 2636 8857 2670 8891
rect 2973 8857 3007 8891
rect 3341 8857 3375 8891
rect 5396 8857 5430 8891
rect 1501 8789 1535 8823
rect 7481 8789 7515 8823
rect 8585 8789 8619 8823
rect 5733 8585 5767 8619
rect 6193 8585 6227 8619
rect 2145 8517 2179 8551
rect 4997 8517 5031 8551
rect 5181 8517 5215 8551
rect 1685 8449 1719 8483
rect 1961 8449 1995 8483
rect 2513 8449 2547 8483
rect 2697 8449 2731 8483
rect 2973 8449 3007 8483
rect 3249 8449 3283 8483
rect 3341 8449 3375 8483
rect 3597 8449 3631 8483
rect 5825 8449 5859 8483
rect 6929 8449 6963 8483
rect 7564 8449 7598 8483
rect 5549 8381 5583 8415
rect 7297 8381 7331 8415
rect 5365 8313 5399 8347
rect 2513 8245 2547 8279
rect 4721 8245 4755 8279
rect 6377 8245 6411 8279
rect 8677 8245 8711 8279
rect 5733 8041 5767 8075
rect 7297 8041 7331 8075
rect 7849 8041 7883 8075
rect 4721 7973 4755 8007
rect 5641 7973 5675 8007
rect 7113 7973 7147 8007
rect 7665 7973 7699 8007
rect 8217 7973 8251 8007
rect 2789 7905 2823 7939
rect 3433 7905 3467 7939
rect 3525 7905 3559 7939
rect 6377 7905 6411 7939
rect 7481 7905 7515 7939
rect 3065 7837 3099 7871
rect 3157 7837 3191 7871
rect 3985 7837 4019 7871
rect 4261 7837 4295 7871
rect 4353 7837 4387 7871
rect 4537 7837 4571 7871
rect 4629 7837 4663 7871
rect 5273 7837 5307 7871
rect 5917 7837 5951 7871
rect 6469 7837 6503 7871
rect 6653 7837 6687 7871
rect 6929 7837 6963 7871
rect 7113 7837 7147 7871
rect 7389 7837 7423 7871
rect 7757 7837 7791 7871
rect 8125 7837 8159 7871
rect 8493 7837 8527 7871
rect 2522 7769 2556 7803
rect 4169 7769 4203 7803
rect 6009 7769 6043 7803
rect 6102 7769 6136 7803
rect 6239 7769 6273 7803
rect 6561 7769 6595 7803
rect 7481 7769 7515 7803
rect 7849 7769 7883 7803
rect 8217 7769 8251 7803
rect 1409 7701 1443 7735
rect 2881 7701 2915 7735
rect 3341 7701 3375 7735
rect 3801 7701 3835 7735
rect 4445 7701 4479 7735
rect 5181 7701 5215 7735
rect 7021 7701 7055 7735
rect 8033 7701 8067 7735
rect 8401 7701 8435 7735
rect 2513 7497 2547 7531
rect 3065 7497 3099 7531
rect 5917 7497 5951 7531
rect 7665 7429 7699 7463
rect 8125 7429 8159 7463
rect 1593 7361 1627 7395
rect 2145 7361 2179 7395
rect 2329 7361 2363 7395
rect 4353 7361 4387 7395
rect 4629 7361 4663 7395
rect 4813 7361 4847 7395
rect 5181 7361 5215 7395
rect 5733 7361 5767 7395
rect 5825 7361 5859 7395
rect 6654 7361 6688 7395
rect 6837 7361 6871 7395
rect 7021 7361 7055 7395
rect 7389 7361 7423 7395
rect 8309 7361 8343 7395
rect 8401 7361 8435 7395
rect 8493 7361 8527 7395
rect 1869 7293 1903 7327
rect 6101 7293 6135 7327
rect 6561 7293 6595 7327
rect 6745 7293 6779 7327
rect 6377 7225 6411 7259
rect 1409 7157 1443 7191
rect 1777 7157 1811 7191
rect 2053 7157 2087 7191
rect 4537 7157 4571 7191
rect 6009 7157 6043 7191
rect 7757 7157 7791 7191
rect 8033 6953 8067 6987
rect 2789 6885 2823 6919
rect 6101 6817 6135 6851
rect 8401 6817 8435 6851
rect 1409 6749 1443 6783
rect 3617 6749 3651 6783
rect 3985 6749 4019 6783
rect 4077 6749 4111 6783
rect 4537 6749 4571 6783
rect 4629 6749 4663 6783
rect 4997 6749 5031 6783
rect 5549 6749 5583 6783
rect 5733 6749 5767 6783
rect 6193 6749 6227 6783
rect 6469 6749 6503 6783
rect 6929 6749 6963 6783
rect 7205 6749 7239 6783
rect 7573 6749 7607 6783
rect 7757 6749 7791 6783
rect 8677 6749 8711 6783
rect 1676 6681 1710 6715
rect 8033 6681 8067 6715
rect 2973 6613 3007 6647
rect 5457 6613 5491 6647
rect 7297 6613 7331 6647
rect 7481 6613 7515 6647
rect 7849 6613 7883 6647
rect 8493 6613 8527 6647
rect 2513 6409 2547 6443
rect 7113 6409 7147 6443
rect 2145 6341 2179 6375
rect 2237 6341 2271 6375
rect 2697 6341 2731 6375
rect 4445 6341 4479 6375
rect 1593 6273 1627 6307
rect 1961 6273 1995 6307
rect 2329 6273 2363 6307
rect 3249 6273 3283 6307
rect 3525 6273 3559 6307
rect 3801 6273 3835 6307
rect 3985 6273 4019 6307
rect 4169 6273 4203 6307
rect 4353 6273 4387 6307
rect 6377 6273 6411 6307
rect 6653 6273 6687 6307
rect 6929 6273 6963 6307
rect 7297 6273 7331 6307
rect 7553 6273 7587 6307
rect 1869 6205 1903 6239
rect 3157 6205 3191 6239
rect 7205 6205 7239 6239
rect 2973 6137 3007 6171
rect 1409 6069 1443 6103
rect 1777 6069 1811 6103
rect 5733 6069 5767 6103
rect 8677 6069 8711 6103
rect 1593 5865 1627 5899
rect 2237 5865 2271 5899
rect 4997 5865 5031 5899
rect 6101 5865 6135 5899
rect 7021 5865 7055 5899
rect 8033 5865 8067 5899
rect 3801 5797 3835 5831
rect 6929 5797 6963 5831
rect 3341 5729 3375 5763
rect 5089 5729 5123 5763
rect 5549 5729 5583 5763
rect 5733 5729 5767 5763
rect 6745 5729 6779 5763
rect 7757 5729 7791 5763
rect 1777 5661 1811 5695
rect 1961 5661 1995 5695
rect 2053 5661 2087 5695
rect 2421 5661 2455 5695
rect 2605 5661 2639 5695
rect 2697 5661 2731 5695
rect 4077 5661 4111 5695
rect 4261 5661 4295 5695
rect 4629 5661 4663 5695
rect 4905 5661 4939 5695
rect 5181 5661 5215 5695
rect 5825 5661 5859 5695
rect 6377 5661 6411 5695
rect 6561 5661 6595 5695
rect 6929 5661 6963 5695
rect 7297 5661 7331 5695
rect 7665 5661 7699 5695
rect 8585 5661 8619 5695
rect 3893 5593 3927 5627
rect 2789 5525 2823 5559
rect 4721 5525 4755 5559
rect 5365 5525 5399 5559
rect 5917 5525 5951 5559
rect 6653 5525 6687 5559
rect 7389 5525 7423 5559
rect 7481 5525 7515 5559
rect 3157 5321 3191 5355
rect 3709 5321 3743 5355
rect 6837 5321 6871 5355
rect 7389 5321 7423 5355
rect 8585 5321 8619 5355
rect 3249 5253 3283 5287
rect 1676 5185 1710 5219
rect 2881 5185 2915 5219
rect 3341 5185 3375 5219
rect 3709 5185 3743 5219
rect 4721 5185 4755 5219
rect 5089 5185 5123 5219
rect 5549 5185 5583 5219
rect 5641 5185 5675 5219
rect 5825 5185 5859 5219
rect 6009 5185 6043 5219
rect 7113 5185 7147 5219
rect 8401 5185 8435 5219
rect 8677 5185 8711 5219
rect 1409 5117 1443 5151
rect 3065 5117 3099 5151
rect 3525 5117 3559 5151
rect 4077 5117 4111 5151
rect 4353 5117 4387 5151
rect 5733 5117 5767 5151
rect 6377 5117 6411 5151
rect 8125 5117 8159 5151
rect 2973 5049 3007 5083
rect 4997 5049 5031 5083
rect 6653 5049 6687 5083
rect 8401 5049 8435 5083
rect 2789 4981 2823 5015
rect 5365 4981 5399 5015
rect 7573 4981 7607 5015
rect 1869 4777 1903 4811
rect 5181 4777 5215 4811
rect 6469 4777 6503 4811
rect 6745 4777 6779 4811
rect 3433 4709 3467 4743
rect 5549 4709 5583 4743
rect 5733 4709 5767 4743
rect 2329 4641 2363 4675
rect 2513 4641 2547 4675
rect 3249 4641 3283 4675
rect 3617 4641 3651 4675
rect 4353 4641 4387 4675
rect 4721 4641 4755 4675
rect 5825 4641 5859 4675
rect 1593 4573 1627 4607
rect 1869 4573 1903 4607
rect 2053 4573 2087 4607
rect 2237 4573 2271 4607
rect 3341 4573 3375 4607
rect 3985 4573 4019 4607
rect 4077 4573 4111 4607
rect 4169 4573 4203 4607
rect 4537 4573 4571 4607
rect 4813 4573 4847 4607
rect 5641 4573 5675 4607
rect 6101 4573 6135 4607
rect 6285 4573 6319 4607
rect 6469 4573 6503 4607
rect 7021 4573 7055 4607
rect 7205 4573 7239 4607
rect 7481 4573 7515 4607
rect 7665 4573 7699 4607
rect 8309 4573 8343 4607
rect 8677 4573 8711 4607
rect 1777 4505 1811 4539
rect 1961 4505 1995 4539
rect 4445 4505 4479 4539
rect 7113 4505 7147 4539
rect 7323 4505 7357 4539
rect 8585 4505 8619 4539
rect 2145 4437 2179 4471
rect 2605 4437 2639 4471
rect 3341 4437 3375 4471
rect 4261 4437 4295 4471
rect 4997 4437 5031 4471
rect 5181 4437 5215 4471
rect 5917 4437 5951 4471
rect 6009 4437 6043 4471
rect 6837 4437 6871 4471
rect 3341 4233 3375 4267
rect 6193 4233 6227 4267
rect 8585 4233 8619 4267
rect 2329 4165 2363 4199
rect 5825 4165 5859 4199
rect 6055 4131 6089 4165
rect 1501 4097 1535 4131
rect 1685 4097 1719 4131
rect 1961 4097 1995 4131
rect 2140 4087 2174 4121
rect 2237 4097 2271 4131
rect 2513 4097 2547 4131
rect 2605 4097 2639 4131
rect 3249 4097 3283 4131
rect 4169 4097 4203 4131
rect 4997 4097 5031 4131
rect 5089 4097 5123 4131
rect 5457 4097 5491 4131
rect 6377 4097 6411 4131
rect 6561 4097 6595 4131
rect 6653 4097 6687 4131
rect 6745 4097 6779 4131
rect 7021 4097 7055 4131
rect 7277 4097 7311 4131
rect 8677 4097 8711 4131
rect 3985 4029 4019 4063
rect 1685 3961 1719 3995
rect 6929 3961 6963 3995
rect 8401 3961 8435 3995
rect 1869 3893 1903 3927
rect 2513 3893 2547 3927
rect 5641 3893 5675 3927
rect 6009 3893 6043 3927
rect 2881 3689 2915 3723
rect 4353 3689 4387 3723
rect 6837 3689 6871 3723
rect 7205 3689 7239 3723
rect 2789 3621 2823 3655
rect 3341 3621 3375 3655
rect 5181 3621 5215 3655
rect 1409 3553 1443 3587
rect 3065 3553 3099 3587
rect 7297 3553 7331 3587
rect 1676 3485 1710 3519
rect 2881 3485 2915 3519
rect 3157 3485 3191 3519
rect 3249 3485 3283 3519
rect 3617 3485 3651 3519
rect 3801 3485 3835 3519
rect 4169 3485 4203 3519
rect 4261 3485 4295 3519
rect 4537 3485 4571 3519
rect 4629 3485 4663 3519
rect 4721 3485 4755 3519
rect 5089 3485 5123 3519
rect 5365 3485 5399 3519
rect 7021 3485 7055 3519
rect 7205 3485 7239 3519
rect 7553 3485 7587 3519
rect 3341 3417 3375 3451
rect 5632 3417 5666 3451
rect 3525 3349 3559 3383
rect 3893 3349 3927 3383
rect 3985 3349 4019 3383
rect 4077 3349 4111 3383
rect 4997 3349 5031 3383
rect 6745 3349 6779 3383
rect 8677 3349 8711 3383
rect 6837 3145 6871 3179
rect 8033 3145 8067 3179
rect 8217 3145 8251 3179
rect 2605 3077 2639 3111
rect 4353 3077 4387 3111
rect 5181 3077 5215 3111
rect 6469 3077 6503 3111
rect 6699 3043 6733 3077
rect 1795 3009 1829 3043
rect 2053 3009 2087 3043
rect 2329 3009 2363 3043
rect 2513 3009 2547 3043
rect 5365 3009 5399 3043
rect 5457 3009 5491 3043
rect 6929 3009 6963 3043
rect 7205 3009 7239 3043
rect 7573 3009 7607 3043
rect 8309 3009 8343 3043
rect 8401 3009 8435 3043
rect 2421 2941 2455 2975
rect 4997 2941 5031 2975
rect 5641 2941 5675 2975
rect 7941 2941 7975 2975
rect 8585 2873 8619 2907
rect 1501 2805 1535 2839
rect 2237 2805 2271 2839
rect 4445 2805 4479 2839
rect 5181 2805 5215 2839
rect 6193 2805 6227 2839
rect 6653 2805 6687 2839
rect 7481 2805 7515 2839
rect 1409 2601 1443 2635
rect 3893 2601 3927 2635
rect 6653 2601 6687 2635
rect 7021 2601 7055 2635
rect 2789 2465 2823 2499
rect 3065 2465 3099 2499
rect 6377 2465 6411 2499
rect 8125 2465 8159 2499
rect 2533 2397 2567 2431
rect 2968 2397 3002 2431
rect 3341 2397 3375 2431
rect 3433 2397 3467 2431
rect 3617 2397 3651 2431
rect 5273 2397 5307 2431
rect 5549 2397 5583 2431
rect 5733 2397 5767 2431
rect 5825 2397 5859 2431
rect 5917 2397 5951 2431
rect 6745 2397 6779 2431
rect 6929 2397 6963 2431
rect 7205 2397 7239 2431
rect 7389 2397 7423 2431
rect 7665 2397 7699 2431
rect 7757 2397 7791 2431
rect 7941 2397 7975 2431
rect 8217 2397 8251 2431
rect 8309 2397 8343 2431
rect 8401 2397 8435 2431
rect 3065 2329 3099 2363
rect 3157 2329 3191 2363
rect 5028 2329 5062 2363
rect 6193 2329 6227 2363
rect 8493 2329 8527 2363
rect 3525 2261 3559 2295
rect 6469 2261 6503 2295
rect 7481 2261 7515 2295
rect 8033 2261 8067 2295
<< metal1 >>
rect 1104 9818 9016 9840
rect 1104 9766 2599 9818
rect 2651 9766 2663 9818
rect 2715 9766 2727 9818
rect 2779 9766 2791 9818
rect 2843 9766 2855 9818
rect 2907 9766 4577 9818
rect 4629 9766 4641 9818
rect 4693 9766 4705 9818
rect 4757 9766 4769 9818
rect 4821 9766 4833 9818
rect 4885 9766 6555 9818
rect 6607 9766 6619 9818
rect 6671 9766 6683 9818
rect 6735 9766 6747 9818
rect 6799 9766 6811 9818
rect 6863 9766 8533 9818
rect 8585 9766 8597 9818
rect 8649 9766 8661 9818
rect 8713 9766 8725 9818
rect 8777 9766 8789 9818
rect 8841 9766 9016 9818
rect 1104 9744 9016 9766
rect 2409 9707 2467 9713
rect 2409 9673 2421 9707
rect 2455 9704 2467 9707
rect 2682 9704 2688 9716
rect 2455 9676 2688 9704
rect 2455 9673 2467 9676
rect 2409 9667 2467 9673
rect 2682 9664 2688 9676
rect 2740 9664 2746 9716
rect 5537 9707 5595 9713
rect 5537 9673 5549 9707
rect 5583 9673 5595 9707
rect 5905 9707 5963 9713
rect 5905 9704 5917 9707
rect 5537 9667 5595 9673
rect 5736 9676 5917 9704
rect 2038 9596 2044 9648
rect 2096 9636 2102 9648
rect 3421 9639 3479 9645
rect 3421 9636 3433 9639
rect 2096 9608 3433 9636
rect 2096 9596 2102 9608
rect 3421 9605 3433 9608
rect 3467 9636 3479 9639
rect 5552 9636 5580 9667
rect 3467 9608 5580 9636
rect 3467 9605 3479 9608
rect 3421 9599 3479 9605
rect 1581 9571 1639 9577
rect 1581 9537 1593 9571
rect 1627 9568 1639 9571
rect 1627 9540 3280 9568
rect 1627 9537 1639 9540
rect 1581 9531 1639 9537
rect 1670 9460 1676 9512
rect 1728 9500 1734 9512
rect 1949 9503 2007 9509
rect 1949 9500 1961 9503
rect 1728 9472 1961 9500
rect 1728 9460 1734 9472
rect 1949 9469 1961 9472
rect 1995 9469 2007 9503
rect 1949 9463 2007 9469
rect 1765 9367 1823 9373
rect 1765 9333 1777 9367
rect 1811 9364 1823 9367
rect 1854 9364 1860 9376
rect 1811 9336 1860 9364
rect 1811 9333 1823 9336
rect 1765 9327 1823 9333
rect 1854 9324 1860 9336
rect 1912 9324 1918 9376
rect 1964 9364 1992 9463
rect 2038 9460 2044 9512
rect 2096 9460 2102 9512
rect 2133 9503 2191 9509
rect 2133 9469 2145 9503
rect 2179 9469 2191 9503
rect 2133 9463 2191 9469
rect 2225 9503 2283 9509
rect 2225 9469 2237 9503
rect 2271 9500 2283 9503
rect 2314 9500 2320 9512
rect 2271 9472 2320 9500
rect 2271 9469 2283 9472
rect 2225 9463 2283 9469
rect 2148 9432 2176 9463
rect 2314 9460 2320 9472
rect 2372 9460 2378 9512
rect 2406 9460 2412 9512
rect 2464 9460 2470 9512
rect 2501 9503 2559 9509
rect 2501 9469 2513 9503
rect 2547 9469 2559 9503
rect 3252 9500 3280 9540
rect 3326 9528 3332 9580
rect 3384 9528 3390 9580
rect 3605 9571 3663 9577
rect 3605 9537 3617 9571
rect 3651 9568 3663 9571
rect 3694 9568 3700 9580
rect 3651 9540 3700 9568
rect 3651 9537 3663 9540
rect 3605 9531 3663 9537
rect 3694 9528 3700 9540
rect 3752 9528 3758 9580
rect 5736 9577 5764 9676
rect 5905 9673 5917 9676
rect 5951 9673 5963 9707
rect 5905 9667 5963 9673
rect 5810 9596 5816 9648
rect 5868 9636 5874 9648
rect 5868 9608 6868 9636
rect 5868 9596 5874 9608
rect 4525 9571 4583 9577
rect 4525 9568 4537 9571
rect 4065 9551 4123 9557
rect 4065 9517 4077 9551
rect 4111 9517 4123 9551
rect 3878 9500 3884 9512
rect 3252 9472 3884 9500
rect 2501 9463 2559 9469
rect 2424 9432 2452 9460
rect 2148 9404 2452 9432
rect 2516 9364 2544 9463
rect 3878 9460 3884 9472
rect 3936 9460 3942 9512
rect 4065 9511 4123 9517
rect 4172 9540 4537 9568
rect 4172 9512 4200 9540
rect 4525 9537 4537 9540
rect 4571 9537 4583 9571
rect 4525 9531 4583 9537
rect 5721 9571 5779 9577
rect 5721 9537 5733 9571
rect 5767 9537 5779 9571
rect 5721 9531 5779 9537
rect 6089 9571 6147 9577
rect 6089 9537 6101 9571
rect 6135 9537 6147 9571
rect 6089 9531 6147 9537
rect 3973 9503 4031 9509
rect 3973 9469 3985 9503
rect 4019 9469 4031 9503
rect 3973 9463 4031 9469
rect 3145 9435 3203 9441
rect 3145 9401 3157 9435
rect 3191 9432 3203 9435
rect 3510 9432 3516 9444
rect 3191 9404 3516 9432
rect 3191 9401 3203 9404
rect 3145 9395 3203 9401
rect 3510 9392 3516 9404
rect 3568 9392 3574 9444
rect 3605 9435 3663 9441
rect 3605 9401 3617 9435
rect 3651 9432 3663 9435
rect 3988 9432 4016 9463
rect 3651 9404 4016 9432
rect 4080 9432 4108 9511
rect 4154 9460 4160 9512
rect 4212 9460 4218 9512
rect 4338 9460 4344 9512
rect 4396 9460 4402 9512
rect 4430 9460 4436 9512
rect 4488 9460 4494 9512
rect 4540 9500 4568 9531
rect 5810 9500 5816 9512
rect 4540 9472 5816 9500
rect 5810 9460 5816 9472
rect 5868 9500 5874 9512
rect 6104 9500 6132 9531
rect 6454 9528 6460 9580
rect 6512 9528 6518 9580
rect 6840 9577 6868 9608
rect 6549 9571 6607 9577
rect 6549 9537 6561 9571
rect 6595 9537 6607 9571
rect 6549 9531 6607 9537
rect 6825 9571 6883 9577
rect 6825 9537 6837 9571
rect 6871 9537 6883 9571
rect 7374 9568 7380 9580
rect 6825 9531 6883 9537
rect 7300 9540 7380 9568
rect 5868 9472 6132 9500
rect 5868 9460 5874 9472
rect 6362 9460 6368 9512
rect 6420 9500 6426 9512
rect 6564 9500 6592 9531
rect 6420 9472 6592 9500
rect 6733 9503 6791 9509
rect 6420 9460 6426 9472
rect 6733 9469 6745 9503
rect 6779 9500 6791 9503
rect 6914 9500 6920 9512
rect 6779 9472 6920 9500
rect 6779 9469 6791 9472
rect 6733 9463 6791 9469
rect 6914 9460 6920 9472
rect 6972 9460 6978 9512
rect 7300 9509 7328 9540
rect 7374 9528 7380 9540
rect 7432 9528 7438 9580
rect 7558 9577 7564 9580
rect 7552 9531 7564 9577
rect 7558 9528 7564 9531
rect 7616 9528 7622 9580
rect 7285 9503 7343 9509
rect 7285 9469 7297 9503
rect 7331 9469 7343 9503
rect 7285 9463 7343 9469
rect 5166 9432 5172 9444
rect 4080 9404 5172 9432
rect 3651 9401 3663 9404
rect 3605 9395 3663 9401
rect 5166 9392 5172 9404
rect 5224 9392 5230 9444
rect 1964 9336 2544 9364
rect 2682 9324 2688 9376
rect 2740 9364 2746 9376
rect 3234 9364 3240 9376
rect 2740 9336 3240 9364
rect 2740 9324 2746 9336
rect 3234 9324 3240 9336
rect 3292 9324 3298 9376
rect 3418 9324 3424 9376
rect 3476 9364 3482 9376
rect 3789 9367 3847 9373
rect 3789 9364 3801 9367
rect 3476 9336 3801 9364
rect 3476 9324 3482 9336
rect 3789 9333 3801 9336
rect 3835 9333 3847 9367
rect 3789 9327 3847 9333
rect 4709 9367 4767 9373
rect 4709 9333 4721 9367
rect 4755 9364 4767 9367
rect 6270 9364 6276 9376
rect 4755 9336 6276 9364
rect 4755 9333 4767 9336
rect 4709 9327 4767 9333
rect 6270 9324 6276 9336
rect 6328 9324 6334 9376
rect 7009 9367 7067 9373
rect 7009 9333 7021 9367
rect 7055 9364 7067 9367
rect 7098 9364 7104 9376
rect 7055 9336 7104 9364
rect 7055 9333 7067 9336
rect 7009 9327 7067 9333
rect 7098 9324 7104 9336
rect 7156 9324 7162 9376
rect 8386 9324 8392 9376
rect 8444 9364 8450 9376
rect 8665 9367 8723 9373
rect 8665 9364 8677 9367
rect 8444 9336 8677 9364
rect 8444 9324 8450 9336
rect 8665 9333 8677 9336
rect 8711 9333 8723 9367
rect 8665 9327 8723 9333
rect 1104 9274 9016 9296
rect 1104 9222 1939 9274
rect 1991 9222 2003 9274
rect 2055 9222 2067 9274
rect 2119 9222 2131 9274
rect 2183 9222 2195 9274
rect 2247 9222 3917 9274
rect 3969 9222 3981 9274
rect 4033 9222 4045 9274
rect 4097 9222 4109 9274
rect 4161 9222 4173 9274
rect 4225 9222 5895 9274
rect 5947 9222 5959 9274
rect 6011 9222 6023 9274
rect 6075 9222 6087 9274
rect 6139 9222 6151 9274
rect 6203 9222 7873 9274
rect 7925 9222 7937 9274
rect 7989 9222 8001 9274
rect 8053 9222 8065 9274
rect 8117 9222 8129 9274
rect 8181 9222 9016 9274
rect 1104 9200 9016 9222
rect 2498 9120 2504 9172
rect 2556 9160 2562 9172
rect 3326 9160 3332 9172
rect 2556 9132 3332 9160
rect 2556 9120 2562 9132
rect 3326 9120 3332 9132
rect 3384 9120 3390 9172
rect 5810 9120 5816 9172
rect 5868 9120 5874 9172
rect 3344 9092 3372 9120
rect 4249 9095 4307 9101
rect 4249 9092 4261 9095
rect 3344 9064 4261 9092
rect 4249 9061 4261 9064
rect 4295 9061 4307 9095
rect 4249 9055 4307 9061
rect 2869 9027 2927 9033
rect 2869 8993 2881 9027
rect 2915 9024 2927 9027
rect 5629 9027 5687 9033
rect 2915 8996 4108 9024
rect 2915 8993 2927 8996
rect 2869 8987 2927 8993
rect 4080 8968 4108 8996
rect 5629 8993 5641 9027
rect 5675 9024 5687 9027
rect 5675 8996 7420 9024
rect 5675 8993 5687 8996
rect 5629 8987 5687 8993
rect 3142 8916 3148 8968
rect 3200 8916 3206 8968
rect 3234 8916 3240 8968
rect 3292 8916 3298 8968
rect 3510 8965 3516 8968
rect 3467 8959 3516 8965
rect 3467 8925 3479 8959
rect 3513 8925 3516 8959
rect 3467 8919 3516 8925
rect 3510 8916 3516 8919
rect 3568 8916 3574 8968
rect 3605 8959 3663 8965
rect 3605 8925 3617 8959
rect 3651 8925 3663 8959
rect 3605 8919 3663 8925
rect 2624 8891 2682 8897
rect 2624 8857 2636 8891
rect 2670 8888 2682 8891
rect 2961 8891 3019 8897
rect 2961 8888 2973 8891
rect 2670 8860 2973 8888
rect 2670 8857 2682 8860
rect 2624 8851 2682 8857
rect 2961 8857 2973 8860
rect 3007 8857 3019 8891
rect 2961 8851 3019 8857
rect 3329 8891 3387 8897
rect 3329 8857 3341 8891
rect 3375 8857 3387 8891
rect 3620 8888 3648 8919
rect 4062 8916 4068 8968
rect 4120 8956 4126 8968
rect 5644 8956 5672 8987
rect 7392 8968 7420 8996
rect 4120 8928 5672 8956
rect 7101 8959 7159 8965
rect 4120 8916 4126 8928
rect 7101 8925 7113 8959
rect 7147 8956 7159 8959
rect 7147 8928 7328 8956
rect 7147 8925 7159 8928
rect 7101 8919 7159 8925
rect 4338 8888 4344 8900
rect 3620 8860 4344 8888
rect 3329 8851 3387 8857
rect 1489 8823 1547 8829
rect 1489 8789 1501 8823
rect 1535 8820 1547 8823
rect 1670 8820 1676 8832
rect 1535 8792 1676 8820
rect 1535 8789 1547 8792
rect 1489 8783 1547 8789
rect 1670 8780 1676 8792
rect 1728 8780 1734 8832
rect 3344 8820 3372 8851
rect 4338 8848 4344 8860
rect 4396 8888 4402 8900
rect 5384 8891 5442 8897
rect 4396 8860 5304 8888
rect 4396 8848 4402 8860
rect 5276 8832 5304 8860
rect 5384 8857 5396 8891
rect 5430 8888 5442 8891
rect 5718 8888 5724 8900
rect 5430 8860 5724 8888
rect 5430 8857 5442 8860
rect 5384 8851 5442 8857
rect 5718 8848 5724 8860
rect 5776 8848 5782 8900
rect 7300 8888 7328 8928
rect 7374 8916 7380 8968
rect 7432 8916 7438 8968
rect 7650 8916 7656 8968
rect 7708 8916 7714 8968
rect 7837 8959 7895 8965
rect 7837 8925 7849 8959
rect 7883 8956 7895 8959
rect 8294 8956 8300 8968
rect 7883 8928 8300 8956
rect 7883 8925 7895 8928
rect 7837 8919 7895 8925
rect 8294 8916 8300 8928
rect 8352 8916 8358 8968
rect 8389 8959 8447 8965
rect 8389 8925 8401 8959
rect 8435 8956 8447 8959
rect 8481 8959 8539 8965
rect 8481 8956 8493 8959
rect 8435 8928 8493 8956
rect 8435 8925 8447 8928
rect 8389 8919 8447 8925
rect 8481 8925 8493 8928
rect 8527 8925 8539 8959
rect 8481 8919 8539 8925
rect 7300 8860 7512 8888
rect 4246 8820 4252 8832
rect 3344 8792 4252 8820
rect 4246 8780 4252 8792
rect 4304 8780 4310 8832
rect 5258 8780 5264 8832
rect 5316 8780 5322 8832
rect 7484 8829 7512 8860
rect 7469 8823 7527 8829
rect 7469 8789 7481 8823
rect 7515 8789 7527 8823
rect 7469 8783 7527 8789
rect 7742 8780 7748 8832
rect 7800 8820 7806 8832
rect 8573 8823 8631 8829
rect 8573 8820 8585 8823
rect 7800 8792 8585 8820
rect 7800 8780 7806 8792
rect 8573 8789 8585 8792
rect 8619 8789 8631 8823
rect 8573 8783 8631 8789
rect 1104 8730 9016 8752
rect 1104 8678 2599 8730
rect 2651 8678 2663 8730
rect 2715 8678 2727 8730
rect 2779 8678 2791 8730
rect 2843 8678 2855 8730
rect 2907 8678 4577 8730
rect 4629 8678 4641 8730
rect 4693 8678 4705 8730
rect 4757 8678 4769 8730
rect 4821 8678 4833 8730
rect 4885 8678 6555 8730
rect 6607 8678 6619 8730
rect 6671 8678 6683 8730
rect 6735 8678 6747 8730
rect 6799 8678 6811 8730
rect 6863 8678 8533 8730
rect 8585 8678 8597 8730
rect 8649 8678 8661 8730
rect 8713 8678 8725 8730
rect 8777 8678 8789 8730
rect 8841 8678 9016 8730
rect 1104 8656 9016 8678
rect 2222 8576 2228 8628
rect 2280 8616 2286 8628
rect 3142 8616 3148 8628
rect 2280 8588 3148 8616
rect 2280 8576 2286 8588
rect 3142 8576 3148 8588
rect 3200 8576 3206 8628
rect 3326 8616 3332 8628
rect 3252 8588 3332 8616
rect 2133 8551 2191 8557
rect 2133 8517 2145 8551
rect 2179 8548 2191 8551
rect 3050 8548 3056 8560
rect 2179 8520 3056 8548
rect 2179 8517 2191 8520
rect 2133 8511 2191 8517
rect 3050 8508 3056 8520
rect 3108 8508 3114 8560
rect 3252 8548 3280 8588
rect 3326 8576 3332 8588
rect 3384 8616 3390 8628
rect 3384 8588 5028 8616
rect 3384 8576 3390 8588
rect 5000 8557 5028 8588
rect 5350 8576 5356 8628
rect 5408 8616 5414 8628
rect 5721 8619 5779 8625
rect 5721 8616 5733 8619
rect 5408 8588 5733 8616
rect 5408 8576 5414 8588
rect 5721 8585 5733 8588
rect 5767 8585 5779 8619
rect 5721 8579 5779 8585
rect 5810 8576 5816 8628
rect 5868 8576 5874 8628
rect 6181 8619 6239 8625
rect 6181 8585 6193 8619
rect 6227 8616 6239 8619
rect 7650 8616 7656 8628
rect 6227 8588 7656 8616
rect 6227 8585 6239 8588
rect 6181 8579 6239 8585
rect 7650 8576 7656 8588
rect 7708 8576 7714 8628
rect 4985 8551 5043 8557
rect 3160 8520 3280 8548
rect 3344 8520 4108 8548
rect 3160 8492 3188 8520
rect 3344 8492 3372 8520
rect 4080 8492 4108 8520
rect 4985 8517 4997 8551
rect 5031 8548 5043 8551
rect 5074 8548 5080 8560
rect 5031 8520 5080 8548
rect 5031 8517 5043 8520
rect 4985 8511 5043 8517
rect 5074 8508 5080 8520
rect 5132 8508 5138 8560
rect 5169 8551 5227 8557
rect 5169 8517 5181 8551
rect 5215 8548 5227 8551
rect 5828 8548 5856 8576
rect 6730 8548 6736 8560
rect 5215 8520 6736 8548
rect 5215 8517 5227 8520
rect 5169 8511 5227 8517
rect 1670 8440 1676 8492
rect 1728 8440 1734 8492
rect 1949 8483 2007 8489
rect 1949 8449 1961 8483
rect 1995 8480 2007 8483
rect 2314 8480 2320 8492
rect 1995 8452 2320 8480
rect 1995 8449 2007 8452
rect 1949 8443 2007 8449
rect 2314 8440 2320 8452
rect 2372 8480 2378 8492
rect 2501 8483 2559 8489
rect 2501 8480 2513 8483
rect 2372 8452 2513 8480
rect 2372 8440 2378 8452
rect 2501 8449 2513 8452
rect 2547 8480 2559 8483
rect 2590 8480 2596 8492
rect 2547 8452 2596 8480
rect 2547 8449 2559 8452
rect 2501 8443 2559 8449
rect 2590 8440 2596 8452
rect 2648 8440 2654 8492
rect 2685 8483 2743 8489
rect 2685 8449 2697 8483
rect 2731 8480 2743 8483
rect 2866 8480 2872 8492
rect 2731 8452 2872 8480
rect 2731 8449 2743 8452
rect 2685 8443 2743 8449
rect 1688 8412 1716 8440
rect 2700 8412 2728 8443
rect 2866 8440 2872 8452
rect 2924 8440 2930 8492
rect 2961 8483 3019 8489
rect 2961 8449 2973 8483
rect 3007 8480 3019 8483
rect 3142 8480 3148 8492
rect 3007 8452 3148 8480
rect 3007 8449 3019 8452
rect 2961 8443 3019 8449
rect 3142 8440 3148 8452
rect 3200 8440 3206 8492
rect 3234 8440 3240 8492
rect 3292 8440 3298 8492
rect 3326 8440 3332 8492
rect 3384 8440 3390 8492
rect 3418 8440 3424 8492
rect 3476 8480 3482 8492
rect 3585 8483 3643 8489
rect 3585 8480 3597 8483
rect 3476 8452 3597 8480
rect 3476 8440 3482 8452
rect 3585 8449 3597 8452
rect 3631 8449 3643 8483
rect 3585 8443 3643 8449
rect 4062 8440 4068 8492
rect 4120 8440 4126 8492
rect 5552 8424 5580 8520
rect 6730 8508 6736 8520
rect 6788 8508 6794 8560
rect 5626 8440 5632 8492
rect 5684 8480 5690 8492
rect 5813 8483 5871 8489
rect 5813 8480 5825 8483
rect 5684 8452 5825 8480
rect 5684 8440 5690 8452
rect 5813 8449 5825 8452
rect 5859 8449 5871 8483
rect 5813 8443 5871 8449
rect 6638 8440 6644 8492
rect 6696 8480 6702 8492
rect 7558 8489 7564 8492
rect 6917 8483 6975 8489
rect 6917 8480 6929 8483
rect 6696 8452 6929 8480
rect 6696 8440 6702 8452
rect 6917 8449 6929 8452
rect 6963 8449 6975 8483
rect 7552 8480 7564 8489
rect 7519 8452 7564 8480
rect 6917 8443 6975 8449
rect 7552 8443 7564 8452
rect 7558 8440 7564 8443
rect 7616 8440 7622 8492
rect 1688 8384 2728 8412
rect 5534 8372 5540 8424
rect 5592 8372 5598 8424
rect 7282 8372 7288 8424
rect 7340 8372 7346 8424
rect 5353 8347 5411 8353
rect 5353 8313 5365 8347
rect 5399 8344 5411 8347
rect 5810 8344 5816 8356
rect 5399 8316 5816 8344
rect 5399 8313 5411 8316
rect 5353 8307 5411 8313
rect 5810 8304 5816 8316
rect 5868 8304 5874 8356
rect 6546 8344 6552 8356
rect 6288 8316 6552 8344
rect 1578 8236 1584 8288
rect 1636 8276 1642 8288
rect 2222 8276 2228 8288
rect 1636 8248 2228 8276
rect 1636 8236 1642 8248
rect 2222 8236 2228 8248
rect 2280 8276 2286 8288
rect 2501 8279 2559 8285
rect 2501 8276 2513 8279
rect 2280 8248 2513 8276
rect 2280 8236 2286 8248
rect 2501 8245 2513 8248
rect 2547 8245 2559 8279
rect 2501 8239 2559 8245
rect 2590 8236 2596 8288
rect 2648 8276 2654 8288
rect 3694 8276 3700 8288
rect 2648 8248 3700 8276
rect 2648 8236 2654 8248
rect 3694 8236 3700 8248
rect 3752 8276 3758 8288
rect 4430 8276 4436 8288
rect 3752 8248 4436 8276
rect 3752 8236 3758 8248
rect 4430 8236 4436 8248
rect 4488 8276 4494 8288
rect 4709 8279 4767 8285
rect 4709 8276 4721 8279
rect 4488 8248 4721 8276
rect 4488 8236 4494 8248
rect 4709 8245 4721 8248
rect 4755 8276 4767 8279
rect 5258 8276 5264 8288
rect 4755 8248 5264 8276
rect 4755 8245 4767 8248
rect 4709 8239 4767 8245
rect 5258 8236 5264 8248
rect 5316 8236 5322 8288
rect 5442 8236 5448 8288
rect 5500 8276 5506 8288
rect 6288 8276 6316 8316
rect 6546 8304 6552 8316
rect 6604 8304 6610 8356
rect 5500 8248 6316 8276
rect 5500 8236 5506 8248
rect 6362 8236 6368 8288
rect 6420 8236 6426 8288
rect 7190 8236 7196 8288
rect 7248 8276 7254 8288
rect 8386 8276 8392 8288
rect 7248 8248 8392 8276
rect 7248 8236 7254 8248
rect 8386 8236 8392 8248
rect 8444 8236 8450 8288
rect 8662 8236 8668 8288
rect 8720 8236 8726 8288
rect 1104 8186 9016 8208
rect 1104 8134 1939 8186
rect 1991 8134 2003 8186
rect 2055 8134 2067 8186
rect 2119 8134 2131 8186
rect 2183 8134 2195 8186
rect 2247 8134 3917 8186
rect 3969 8134 3981 8186
rect 4033 8134 4045 8186
rect 4097 8134 4109 8186
rect 4161 8134 4173 8186
rect 4225 8134 5895 8186
rect 5947 8134 5959 8186
rect 6011 8134 6023 8186
rect 6075 8134 6087 8186
rect 6139 8134 6151 8186
rect 6203 8134 7873 8186
rect 7925 8134 7937 8186
rect 7989 8134 8001 8186
rect 8053 8134 8065 8186
rect 8117 8134 8129 8186
rect 8181 8134 9016 8186
rect 1104 8112 9016 8134
rect 3804 8044 5580 8072
rect 2866 7964 2872 8016
rect 2924 8004 2930 8016
rect 2924 7976 3464 8004
rect 2924 7964 2930 7976
rect 2777 7939 2835 7945
rect 2777 7905 2789 7939
rect 2823 7936 2835 7939
rect 3326 7936 3332 7948
rect 2823 7908 3332 7936
rect 2823 7905 2835 7908
rect 2777 7899 2835 7905
rect 3326 7896 3332 7908
rect 3384 7896 3390 7948
rect 3436 7945 3464 7976
rect 3421 7939 3479 7945
rect 3421 7905 3433 7939
rect 3467 7905 3479 7939
rect 3421 7899 3479 7905
rect 3513 7939 3571 7945
rect 3513 7905 3525 7939
rect 3559 7936 3571 7939
rect 3694 7936 3700 7948
rect 3559 7908 3700 7936
rect 3559 7905 3571 7908
rect 3513 7899 3571 7905
rect 3694 7896 3700 7908
rect 3752 7896 3758 7948
rect 3053 7871 3111 7877
rect 3053 7868 3065 7871
rect 2056 7840 3065 7868
rect 2056 7744 2084 7840
rect 3053 7837 3065 7840
rect 3099 7837 3111 7871
rect 3053 7831 3111 7837
rect 3145 7871 3203 7877
rect 3145 7837 3157 7871
rect 3191 7837 3203 7871
rect 3804 7868 3832 8044
rect 5552 8016 5580 8044
rect 5718 8032 5724 8084
rect 5776 8032 5782 8084
rect 6362 8032 6368 8084
rect 6420 8032 6426 8084
rect 6730 8032 6736 8084
rect 6788 8032 6794 8084
rect 7190 8032 7196 8084
rect 7248 8072 7254 8084
rect 7285 8075 7343 8081
rect 7285 8072 7297 8075
rect 7248 8044 7297 8072
rect 7248 8032 7254 8044
rect 7285 8041 7297 8044
rect 7331 8041 7343 8075
rect 7285 8035 7343 8041
rect 7558 8032 7564 8084
rect 7616 8072 7622 8084
rect 7837 8075 7895 8081
rect 7837 8072 7849 8075
rect 7616 8044 7849 8072
rect 7616 8032 7622 8044
rect 7837 8041 7849 8044
rect 7883 8041 7895 8075
rect 7837 8035 7895 8041
rect 3878 7964 3884 8016
rect 3936 8004 3942 8016
rect 4709 8007 4767 8013
rect 4709 8004 4721 8007
rect 3936 7976 4721 8004
rect 3936 7964 3942 7976
rect 4709 7973 4721 7976
rect 4755 7973 4767 8007
rect 4709 7967 4767 7973
rect 5534 7964 5540 8016
rect 5592 8004 5598 8016
rect 5629 8007 5687 8013
rect 5629 8004 5641 8007
rect 5592 7976 5641 8004
rect 5592 7964 5598 7976
rect 5629 7973 5641 7976
rect 5675 7973 5687 8007
rect 6178 8004 6184 8016
rect 5629 7967 5687 7973
rect 5828 7976 6184 8004
rect 4982 7936 4988 7948
rect 4264 7908 4988 7936
rect 4264 7877 4292 7908
rect 4982 7896 4988 7908
rect 5040 7896 5046 7948
rect 5350 7896 5356 7948
rect 5408 7936 5414 7948
rect 5828 7936 5856 7976
rect 6178 7964 6184 7976
rect 6236 7964 6242 8016
rect 6380 7945 6408 8032
rect 6748 8004 6776 8032
rect 6472 7976 6776 8004
rect 7101 8007 7159 8013
rect 6365 7939 6423 7945
rect 5408 7908 5856 7936
rect 5920 7908 6316 7936
rect 5408 7896 5414 7908
rect 3973 7871 4031 7877
rect 3973 7868 3985 7871
rect 3804 7840 3985 7868
rect 3145 7831 3203 7837
rect 3973 7837 3985 7840
rect 4019 7837 4031 7871
rect 3973 7831 4031 7837
rect 4249 7871 4307 7877
rect 4249 7837 4261 7871
rect 4295 7837 4307 7871
rect 4249 7831 4307 7837
rect 4341 7871 4399 7877
rect 4341 7837 4353 7871
rect 4387 7837 4399 7871
rect 4341 7831 4399 7837
rect 2498 7760 2504 7812
rect 2556 7809 2562 7812
rect 2556 7763 2568 7809
rect 3160 7800 3188 7831
rect 4157 7803 4215 7809
rect 4157 7800 4169 7803
rect 2746 7772 3188 7800
rect 3712 7772 4169 7800
rect 2556 7760 2562 7763
rect 1397 7735 1455 7741
rect 1397 7701 1409 7735
rect 1443 7732 1455 7735
rect 2038 7732 2044 7744
rect 1443 7704 2044 7732
rect 1443 7701 1455 7704
rect 1397 7695 1455 7701
rect 2038 7692 2044 7704
rect 2096 7692 2102 7744
rect 2406 7692 2412 7744
rect 2464 7732 2470 7744
rect 2746 7732 2774 7772
rect 3712 7744 3740 7772
rect 4157 7769 4169 7772
rect 4203 7800 4215 7803
rect 4356 7800 4384 7831
rect 4430 7828 4436 7880
rect 4488 7868 4494 7880
rect 4525 7871 4583 7877
rect 4525 7868 4537 7871
rect 4488 7840 4537 7868
rect 4488 7828 4494 7840
rect 4525 7837 4537 7840
rect 4571 7868 4583 7871
rect 4617 7871 4675 7877
rect 4617 7868 4629 7871
rect 4571 7840 4629 7868
rect 4571 7837 4583 7840
rect 4525 7831 4583 7837
rect 4617 7837 4629 7840
rect 4663 7837 4675 7871
rect 4617 7831 4675 7837
rect 5074 7828 5080 7880
rect 5132 7868 5138 7880
rect 5920 7877 5948 7908
rect 5261 7871 5319 7877
rect 5261 7868 5273 7871
rect 5132 7840 5273 7868
rect 5132 7828 5138 7840
rect 5261 7837 5273 7840
rect 5307 7837 5319 7871
rect 5261 7831 5319 7837
rect 5905 7871 5963 7877
rect 5905 7837 5917 7871
rect 5951 7837 5963 7871
rect 6288 7868 6316 7908
rect 6365 7905 6377 7939
rect 6411 7905 6423 7939
rect 6365 7899 6423 7905
rect 6472 7877 6500 7976
rect 7101 7973 7113 8007
rect 7147 7973 7159 8007
rect 7101 7967 7159 7973
rect 6546 7896 6552 7948
rect 6604 7936 6610 7948
rect 7116 7936 7144 7967
rect 7374 7964 7380 8016
rect 7432 8004 7438 8016
rect 7650 8004 7656 8016
rect 7432 7976 7656 8004
rect 7432 7964 7438 7976
rect 7650 7964 7656 7976
rect 7708 7964 7714 8016
rect 7742 7964 7748 8016
rect 7800 8004 7806 8016
rect 8205 8007 8263 8013
rect 7800 7976 7880 8004
rect 7800 7964 7806 7976
rect 7469 7939 7527 7945
rect 7469 7936 7481 7939
rect 6604 7908 6960 7936
rect 7116 7908 7481 7936
rect 6604 7896 6610 7908
rect 6457 7871 6515 7877
rect 6288 7840 6408 7868
rect 5905 7831 5963 7837
rect 4203 7772 4384 7800
rect 4203 7769 4215 7772
rect 4157 7763 4215 7769
rect 5994 7760 6000 7812
rect 6052 7760 6058 7812
rect 6086 7760 6092 7812
rect 6144 7760 6150 7812
rect 6178 7760 6184 7812
rect 6236 7809 6242 7812
rect 6236 7803 6285 7809
rect 6236 7769 6239 7803
rect 6273 7769 6285 7803
rect 6380 7800 6408 7840
rect 6457 7837 6469 7871
rect 6503 7837 6515 7871
rect 6457 7831 6515 7837
rect 6638 7828 6644 7880
rect 6696 7828 6702 7880
rect 6932 7877 6960 7908
rect 7469 7905 7481 7908
rect 7515 7905 7527 7939
rect 7469 7899 7527 7905
rect 7558 7896 7564 7948
rect 7616 7896 7622 7948
rect 6917 7871 6975 7877
rect 6917 7837 6929 7871
rect 6963 7837 6975 7871
rect 6917 7831 6975 7837
rect 7101 7871 7159 7877
rect 7101 7837 7113 7871
rect 7147 7868 7159 7871
rect 7377 7871 7435 7877
rect 7147 7840 7236 7868
rect 7147 7837 7159 7840
rect 7101 7831 7159 7837
rect 6549 7803 6607 7809
rect 6549 7800 6561 7803
rect 6380 7772 6561 7800
rect 6236 7763 6285 7769
rect 6549 7769 6561 7772
rect 6595 7769 6607 7803
rect 6549 7763 6607 7769
rect 6236 7760 6242 7763
rect 2464 7704 2774 7732
rect 2869 7735 2927 7741
rect 2464 7692 2470 7704
rect 2869 7701 2881 7735
rect 2915 7732 2927 7735
rect 2958 7732 2964 7744
rect 2915 7704 2964 7732
rect 2915 7701 2927 7704
rect 2869 7695 2927 7701
rect 2958 7692 2964 7704
rect 3016 7692 3022 7744
rect 3142 7692 3148 7744
rect 3200 7732 3206 7744
rect 3329 7735 3387 7741
rect 3329 7732 3341 7735
rect 3200 7704 3341 7732
rect 3200 7692 3206 7704
rect 3329 7701 3341 7704
rect 3375 7732 3387 7735
rect 3418 7732 3424 7744
rect 3375 7704 3424 7732
rect 3375 7701 3387 7704
rect 3329 7695 3387 7701
rect 3418 7692 3424 7704
rect 3476 7692 3482 7744
rect 3694 7692 3700 7744
rect 3752 7692 3758 7744
rect 3786 7692 3792 7744
rect 3844 7692 3850 7744
rect 4430 7692 4436 7744
rect 4488 7692 4494 7744
rect 5074 7692 5080 7744
rect 5132 7732 5138 7744
rect 5169 7735 5227 7741
rect 5169 7732 5181 7735
rect 5132 7704 5181 7732
rect 5132 7692 5138 7704
rect 5169 7701 5181 7704
rect 5215 7701 5227 7735
rect 5169 7695 5227 7701
rect 6362 7692 6368 7744
rect 6420 7732 6426 7744
rect 6656 7732 6684 7828
rect 6420 7704 6684 7732
rect 6420 7692 6426 7704
rect 7006 7692 7012 7744
rect 7064 7692 7070 7744
rect 7208 7732 7236 7840
rect 7377 7837 7389 7871
rect 7423 7868 7435 7871
rect 7576 7868 7604 7896
rect 7423 7840 7604 7868
rect 7745 7871 7803 7877
rect 7423 7837 7435 7840
rect 7377 7831 7435 7837
rect 7745 7837 7757 7871
rect 7791 7870 7803 7871
rect 7852 7870 7880 7976
rect 8205 7973 8217 8007
rect 8251 7973 8263 8007
rect 8205 7967 8263 7973
rect 8220 7936 8248 7967
rect 7791 7842 7880 7870
rect 7944 7908 8248 7936
rect 7791 7837 7803 7842
rect 7745 7831 7803 7837
rect 7466 7760 7472 7812
rect 7524 7760 7530 7812
rect 7558 7760 7564 7812
rect 7616 7800 7622 7812
rect 7837 7803 7895 7809
rect 7837 7800 7849 7803
rect 7616 7772 7849 7800
rect 7616 7760 7622 7772
rect 7837 7769 7849 7772
rect 7883 7769 7895 7803
rect 7837 7763 7895 7769
rect 7944 7732 7972 7908
rect 8018 7828 8024 7880
rect 8076 7868 8082 7880
rect 8113 7871 8171 7877
rect 8113 7868 8125 7871
rect 8076 7840 8125 7868
rect 8076 7828 8082 7840
rect 8113 7837 8125 7840
rect 8159 7837 8171 7871
rect 8113 7831 8171 7837
rect 8386 7828 8392 7880
rect 8444 7868 8450 7880
rect 8481 7871 8539 7877
rect 8481 7868 8493 7871
rect 8444 7840 8493 7868
rect 8444 7828 8450 7840
rect 8481 7837 8493 7840
rect 8527 7837 8539 7871
rect 8481 7831 8539 7837
rect 8205 7803 8263 7809
rect 8205 7769 8217 7803
rect 8251 7800 8263 7803
rect 8294 7800 8300 7812
rect 8251 7772 8300 7800
rect 8251 7769 8263 7772
rect 8205 7763 8263 7769
rect 8294 7760 8300 7772
rect 8352 7760 8358 7812
rect 7208 7704 7972 7732
rect 8021 7735 8079 7741
rect 8021 7701 8033 7735
rect 8067 7732 8079 7735
rect 8110 7732 8116 7744
rect 8067 7704 8116 7732
rect 8067 7701 8079 7704
rect 8021 7695 8079 7701
rect 8110 7692 8116 7704
rect 8168 7732 8174 7744
rect 8389 7735 8447 7741
rect 8389 7732 8401 7735
rect 8168 7704 8401 7732
rect 8168 7692 8174 7704
rect 8389 7701 8401 7704
rect 8435 7732 8447 7735
rect 8662 7732 8668 7744
rect 8435 7704 8668 7732
rect 8435 7701 8447 7704
rect 8389 7695 8447 7701
rect 8662 7692 8668 7704
rect 8720 7692 8726 7744
rect 1104 7642 9016 7664
rect 1104 7590 2599 7642
rect 2651 7590 2663 7642
rect 2715 7590 2727 7642
rect 2779 7590 2791 7642
rect 2843 7590 2855 7642
rect 2907 7590 4577 7642
rect 4629 7590 4641 7642
rect 4693 7590 4705 7642
rect 4757 7590 4769 7642
rect 4821 7590 4833 7642
rect 4885 7590 6555 7642
rect 6607 7590 6619 7642
rect 6671 7590 6683 7642
rect 6735 7590 6747 7642
rect 6799 7590 6811 7642
rect 6863 7590 8533 7642
rect 8585 7590 8597 7642
rect 8649 7590 8661 7642
rect 8713 7590 8725 7642
rect 8777 7590 8789 7642
rect 8841 7590 9016 7642
rect 1104 7568 9016 7590
rect 2406 7488 2412 7540
rect 2464 7528 2470 7540
rect 2501 7531 2559 7537
rect 2501 7528 2513 7531
rect 2464 7500 2513 7528
rect 2464 7488 2470 7500
rect 2501 7497 2513 7500
rect 2547 7497 2559 7531
rect 2501 7491 2559 7497
rect 2774 7488 2780 7540
rect 2832 7528 2838 7540
rect 3053 7531 3111 7537
rect 3053 7528 3065 7531
rect 2832 7500 3065 7528
rect 2832 7488 2838 7500
rect 3053 7497 3065 7500
rect 3099 7528 3111 7531
rect 3326 7528 3332 7540
rect 3099 7500 3332 7528
rect 3099 7497 3111 7500
rect 3053 7491 3111 7497
rect 3326 7488 3332 7500
rect 3384 7488 3390 7540
rect 3510 7488 3516 7540
rect 3568 7528 3574 7540
rect 4338 7528 4344 7540
rect 3568 7500 4344 7528
rect 3568 7488 3574 7500
rect 4338 7488 4344 7500
rect 4396 7488 4402 7540
rect 5905 7531 5963 7537
rect 5905 7497 5917 7531
rect 5951 7528 5963 7531
rect 7190 7528 7196 7540
rect 5951 7500 7196 7528
rect 5951 7497 5963 7500
rect 5905 7491 5963 7497
rect 7190 7488 7196 7500
rect 7248 7528 7254 7540
rect 7248 7500 7787 7528
rect 7248 7488 7254 7500
rect 1596 7432 3924 7460
rect 1596 7401 1624 7432
rect 1581 7395 1639 7401
rect 1581 7361 1593 7395
rect 1627 7361 1639 7395
rect 1581 7355 1639 7361
rect 2038 7352 2044 7404
rect 2096 7392 2102 7404
rect 2133 7395 2191 7401
rect 2133 7392 2145 7395
rect 2096 7364 2145 7392
rect 2096 7352 2102 7364
rect 2133 7361 2145 7364
rect 2179 7361 2191 7395
rect 2133 7355 2191 7361
rect 2317 7395 2375 7401
rect 2317 7361 2329 7395
rect 2363 7392 2375 7395
rect 3234 7392 3240 7404
rect 2363 7364 3240 7392
rect 2363 7361 2375 7364
rect 2317 7355 2375 7361
rect 1857 7327 1915 7333
rect 1857 7293 1869 7327
rect 1903 7324 1915 7327
rect 2148 7324 2176 7355
rect 3234 7352 3240 7364
rect 3292 7392 3298 7404
rect 3786 7392 3792 7404
rect 3292 7364 3792 7392
rect 3292 7352 3298 7364
rect 3786 7352 3792 7364
rect 3844 7352 3850 7404
rect 2406 7324 2412 7336
rect 1903 7296 2084 7324
rect 2148 7296 2412 7324
rect 1903 7293 1915 7296
rect 1857 7287 1915 7293
rect 1394 7148 1400 7200
rect 1452 7148 1458 7200
rect 1578 7148 1584 7200
rect 1636 7188 1642 7200
rect 2056 7197 2084 7296
rect 2406 7284 2412 7296
rect 2464 7284 2470 7336
rect 3896 7256 3924 7432
rect 5258 7420 5264 7472
rect 5316 7460 5322 7472
rect 5316 7432 6224 7460
rect 5316 7420 5322 7432
rect 4338 7352 4344 7404
rect 4396 7352 4402 7404
rect 4614 7352 4620 7404
rect 4672 7352 4678 7404
rect 4801 7395 4859 7401
rect 4801 7361 4813 7395
rect 4847 7361 4859 7395
rect 4801 7355 4859 7361
rect 4246 7284 4252 7336
rect 4304 7284 4310 7336
rect 4522 7284 4528 7336
rect 4580 7324 4586 7336
rect 4816 7324 4844 7355
rect 4890 7352 4896 7404
rect 4948 7392 4954 7404
rect 5169 7395 5227 7401
rect 5169 7392 5181 7395
rect 4948 7364 5181 7392
rect 4948 7352 4954 7364
rect 5169 7361 5181 7364
rect 5215 7361 5227 7395
rect 5721 7395 5779 7401
rect 5721 7392 5733 7395
rect 5169 7355 5227 7361
rect 5460 7364 5733 7392
rect 5460 7336 5488 7364
rect 5721 7361 5733 7364
rect 5767 7361 5779 7395
rect 5721 7355 5779 7361
rect 5813 7395 5871 7401
rect 5813 7361 5825 7395
rect 5859 7392 5871 7395
rect 5902 7392 5908 7404
rect 5859 7364 5908 7392
rect 5859 7361 5871 7364
rect 5813 7355 5871 7361
rect 5902 7352 5908 7364
rect 5960 7352 5966 7404
rect 4580 7296 4844 7324
rect 4580 7284 4586 7296
rect 5258 7284 5264 7336
rect 5316 7284 5322 7336
rect 5442 7284 5448 7336
rect 5500 7284 5506 7336
rect 5534 7284 5540 7336
rect 5592 7324 5598 7336
rect 6089 7327 6147 7333
rect 6089 7324 6101 7327
rect 5592 7296 6101 7324
rect 5592 7284 5598 7296
rect 6089 7293 6101 7296
rect 6135 7293 6147 7327
rect 6196 7324 6224 7432
rect 7098 7420 7104 7472
rect 7156 7460 7162 7472
rect 7466 7460 7472 7472
rect 7156 7432 7472 7460
rect 7156 7420 7162 7432
rect 7466 7420 7472 7432
rect 7524 7460 7530 7472
rect 7653 7463 7711 7469
rect 7653 7460 7665 7463
rect 7524 7432 7665 7460
rect 7524 7420 7530 7432
rect 7653 7429 7665 7432
rect 7699 7429 7711 7463
rect 7759 7460 7787 7500
rect 7834 7488 7840 7540
rect 7892 7528 7898 7540
rect 8294 7528 8300 7540
rect 7892 7500 8300 7528
rect 7892 7488 7898 7500
rect 8294 7488 8300 7500
rect 8352 7488 8358 7540
rect 8113 7463 8171 7469
rect 8113 7460 8125 7463
rect 7759 7432 8125 7460
rect 7653 7423 7711 7429
rect 8113 7429 8125 7432
rect 8159 7429 8171 7463
rect 8113 7423 8171 7429
rect 8202 7420 8208 7472
rect 8260 7460 8266 7472
rect 8260 7432 8432 7460
rect 8260 7420 8266 7432
rect 6362 7352 6368 7404
rect 6420 7392 6426 7404
rect 6642 7398 6700 7401
rect 6564 7395 6700 7398
rect 6564 7392 6654 7395
rect 6420 7370 6654 7392
rect 6420 7364 6592 7370
rect 6420 7352 6426 7364
rect 6642 7361 6654 7370
rect 6688 7361 6700 7395
rect 6642 7355 6700 7361
rect 6822 7352 6828 7404
rect 6880 7392 6886 7404
rect 7009 7395 7067 7401
rect 7009 7392 7021 7395
rect 6880 7364 7021 7392
rect 6880 7352 6886 7364
rect 7009 7361 7021 7364
rect 7055 7361 7067 7395
rect 7009 7355 7067 7361
rect 7377 7395 7435 7401
rect 7377 7361 7389 7395
rect 7423 7392 7435 7395
rect 7423 7364 7972 7392
rect 7423 7361 7435 7364
rect 7377 7355 7435 7361
rect 6549 7327 6607 7333
rect 6549 7324 6561 7327
rect 6196 7296 6561 7324
rect 6089 7287 6147 7293
rect 6549 7293 6561 7296
rect 6595 7293 6607 7327
rect 6549 7287 6607 7293
rect 6730 7284 6736 7336
rect 6788 7284 6794 7336
rect 4264 7256 4292 7284
rect 5276 7256 5304 7284
rect 5552 7256 5580 7284
rect 6365 7259 6423 7265
rect 6365 7256 6377 7259
rect 3896 7228 5580 7256
rect 5635 7228 6377 7256
rect 1765 7191 1823 7197
rect 1765 7188 1777 7191
rect 1636 7160 1777 7188
rect 1636 7148 1642 7160
rect 1765 7157 1777 7160
rect 1811 7157 1823 7191
rect 1765 7151 1823 7157
rect 2041 7191 2099 7197
rect 2041 7157 2053 7191
rect 2087 7188 2099 7191
rect 3234 7188 3240 7200
rect 2087 7160 3240 7188
rect 2087 7157 2099 7160
rect 2041 7151 2099 7157
rect 3234 7148 3240 7160
rect 3292 7148 3298 7200
rect 4246 7148 4252 7200
rect 4304 7188 4310 7200
rect 4525 7191 4583 7197
rect 4525 7188 4537 7191
rect 4304 7160 4537 7188
rect 4304 7148 4310 7160
rect 4525 7157 4537 7160
rect 4571 7157 4583 7191
rect 4525 7151 4583 7157
rect 5166 7148 5172 7200
rect 5224 7188 5230 7200
rect 5635 7188 5663 7228
rect 6365 7225 6377 7228
rect 6411 7225 6423 7259
rect 7834 7256 7840 7268
rect 6365 7219 6423 7225
rect 6656 7228 7840 7256
rect 5224 7160 5663 7188
rect 5997 7191 6055 7197
rect 5224 7148 5230 7160
rect 5997 7157 6009 7191
rect 6043 7188 6055 7191
rect 6270 7188 6276 7200
rect 6043 7160 6276 7188
rect 6043 7157 6055 7160
rect 5997 7151 6055 7157
rect 6270 7148 6276 7160
rect 6328 7188 6334 7200
rect 6656 7188 6684 7228
rect 7834 7216 7840 7228
rect 7892 7216 7898 7268
rect 6328 7160 6684 7188
rect 6328 7148 6334 7160
rect 7742 7148 7748 7200
rect 7800 7148 7806 7200
rect 7944 7188 7972 7364
rect 8294 7352 8300 7404
rect 8352 7352 8358 7404
rect 8404 7401 8432 7432
rect 8389 7395 8447 7401
rect 8389 7361 8401 7395
rect 8435 7361 8447 7395
rect 8389 7355 8447 7361
rect 8481 7395 8539 7401
rect 8481 7361 8493 7395
rect 8527 7361 8539 7395
rect 8481 7355 8539 7361
rect 8496 7324 8524 7355
rect 8404 7296 8524 7324
rect 8404 7268 8432 7296
rect 8386 7216 8392 7268
rect 8444 7216 8450 7268
rect 8478 7188 8484 7200
rect 7944 7160 8484 7188
rect 8478 7148 8484 7160
rect 8536 7148 8542 7200
rect 1104 7098 9016 7120
rect 1104 7046 1939 7098
rect 1991 7046 2003 7098
rect 2055 7046 2067 7098
rect 2119 7046 2131 7098
rect 2183 7046 2195 7098
rect 2247 7046 3917 7098
rect 3969 7046 3981 7098
rect 4033 7046 4045 7098
rect 4097 7046 4109 7098
rect 4161 7046 4173 7098
rect 4225 7046 5895 7098
rect 5947 7046 5959 7098
rect 6011 7046 6023 7098
rect 6075 7046 6087 7098
rect 6139 7046 6151 7098
rect 6203 7046 7873 7098
rect 7925 7046 7937 7098
rect 7989 7046 8001 7098
rect 8053 7046 8065 7098
rect 8117 7046 8129 7098
rect 8181 7046 9016 7098
rect 1104 7024 9016 7046
rect 6362 6944 6368 6996
rect 6420 6984 6426 6996
rect 6730 6984 6736 6996
rect 6420 6956 6736 6984
rect 6420 6944 6426 6956
rect 6730 6944 6736 6956
rect 6788 6944 6794 6996
rect 8021 6987 8079 6993
rect 8021 6953 8033 6987
rect 8067 6984 8079 6987
rect 8386 6984 8392 6996
rect 8067 6956 8392 6984
rect 8067 6953 8079 6956
rect 8021 6947 8079 6953
rect 8386 6944 8392 6956
rect 8444 6944 8450 6996
rect 2777 6919 2835 6925
rect 2777 6885 2789 6919
rect 2823 6916 2835 6919
rect 2823 6888 3096 6916
rect 2823 6885 2835 6888
rect 2777 6879 2835 6885
rect 1397 6783 1455 6789
rect 1397 6749 1409 6783
rect 1443 6780 1455 6783
rect 2774 6780 2780 6792
rect 1443 6752 2780 6780
rect 1443 6749 1455 6752
rect 1397 6743 1455 6749
rect 2774 6740 2780 6752
rect 2832 6740 2838 6792
rect 1670 6721 1676 6724
rect 1664 6675 1676 6721
rect 1670 6672 1676 6675
rect 1728 6672 1734 6724
rect 3068 6712 3096 6888
rect 3234 6876 3240 6928
rect 3292 6916 3298 6928
rect 3878 6916 3884 6928
rect 3292 6888 3884 6916
rect 3292 6876 3298 6888
rect 3878 6876 3884 6888
rect 3936 6916 3942 6928
rect 4522 6916 4528 6928
rect 3936 6888 4528 6916
rect 3936 6876 3942 6888
rect 4522 6876 4528 6888
rect 4580 6876 4586 6928
rect 5534 6876 5540 6928
rect 5592 6916 5598 6928
rect 5718 6916 5724 6928
rect 5592 6888 5724 6916
rect 5592 6876 5598 6888
rect 5718 6876 5724 6888
rect 5776 6876 5782 6928
rect 5810 6876 5816 6928
rect 5868 6916 5874 6928
rect 6454 6916 6460 6928
rect 5868 6888 6460 6916
rect 5868 6876 5874 6888
rect 6454 6876 6460 6888
rect 6512 6876 6518 6928
rect 4890 6848 4896 6860
rect 3160 6820 4896 6848
rect 3160 6792 3188 6820
rect 4890 6808 4896 6820
rect 4948 6848 4954 6860
rect 6089 6851 6147 6857
rect 4948 6820 5028 6848
rect 4948 6808 4954 6820
rect 3142 6740 3148 6792
rect 3200 6740 3206 6792
rect 3605 6783 3663 6789
rect 3605 6749 3617 6783
rect 3651 6749 3663 6783
rect 3605 6743 3663 6749
rect 3510 6712 3516 6724
rect 3068 6684 3516 6712
rect 3510 6672 3516 6684
rect 3568 6712 3574 6724
rect 3620 6712 3648 6743
rect 3970 6740 3976 6792
rect 4028 6740 4034 6792
rect 4062 6740 4068 6792
rect 4120 6740 4126 6792
rect 4522 6740 4528 6792
rect 4580 6740 4586 6792
rect 4614 6740 4620 6792
rect 4672 6740 4678 6792
rect 5000 6789 5028 6820
rect 5092 6820 5856 6848
rect 4985 6783 5043 6789
rect 4985 6749 4997 6783
rect 5031 6749 5043 6783
rect 4985 6743 5043 6749
rect 4632 6712 4660 6740
rect 3568 6684 4660 6712
rect 3568 6672 3574 6684
rect 1854 6604 1860 6656
rect 1912 6644 1918 6656
rect 2961 6647 3019 6653
rect 2961 6644 2973 6647
rect 1912 6616 2973 6644
rect 1912 6604 1918 6616
rect 2961 6613 2973 6616
rect 3007 6613 3019 6647
rect 2961 6607 3019 6613
rect 4062 6604 4068 6656
rect 4120 6644 4126 6656
rect 5092 6644 5120 6820
rect 5537 6783 5595 6789
rect 5537 6749 5549 6783
rect 5583 6749 5595 6783
rect 5537 6743 5595 6749
rect 5552 6712 5580 6743
rect 5718 6740 5724 6792
rect 5776 6740 5782 6792
rect 5828 6780 5856 6820
rect 6089 6817 6101 6851
rect 6135 6848 6147 6851
rect 7466 6848 7472 6860
rect 6135 6820 7052 6848
rect 6135 6817 6147 6820
rect 6089 6811 6147 6817
rect 7024 6792 7052 6820
rect 7300 6820 7472 6848
rect 6178 6780 6184 6792
rect 5828 6752 6184 6780
rect 6178 6740 6184 6752
rect 6236 6740 6242 6792
rect 6454 6740 6460 6792
rect 6512 6740 6518 6792
rect 6914 6740 6920 6792
rect 6972 6740 6978 6792
rect 7006 6740 7012 6792
rect 7064 6780 7070 6792
rect 7193 6783 7251 6789
rect 7193 6780 7205 6783
rect 7064 6752 7205 6780
rect 7064 6740 7070 6752
rect 7193 6749 7205 6752
rect 7239 6749 7251 6783
rect 7193 6743 7251 6749
rect 7300 6712 7328 6820
rect 7466 6808 7472 6820
rect 7524 6808 7530 6860
rect 8294 6808 8300 6860
rect 8352 6848 8358 6860
rect 8389 6851 8447 6857
rect 8389 6848 8401 6851
rect 8352 6820 8401 6848
rect 8352 6808 8358 6820
rect 8389 6817 8401 6820
rect 8435 6848 8447 6851
rect 8938 6848 8944 6860
rect 8435 6820 8944 6848
rect 8435 6817 8447 6820
rect 8389 6811 8447 6817
rect 8938 6808 8944 6820
rect 8996 6808 9002 6860
rect 7374 6740 7380 6792
rect 7432 6780 7438 6792
rect 7561 6783 7619 6789
rect 7561 6780 7573 6783
rect 7432 6752 7573 6780
rect 7432 6740 7438 6752
rect 7561 6749 7573 6752
rect 7607 6749 7619 6783
rect 7561 6743 7619 6749
rect 7745 6783 7803 6789
rect 7745 6749 7757 6783
rect 7791 6780 7803 6783
rect 8202 6780 8208 6792
rect 7791 6752 8208 6780
rect 7791 6749 7803 6752
rect 7745 6743 7803 6749
rect 8202 6740 8208 6752
rect 8260 6740 8266 6792
rect 8665 6783 8723 6789
rect 8665 6749 8677 6783
rect 8711 6780 8723 6783
rect 9030 6780 9036 6792
rect 8711 6752 9036 6780
rect 8711 6749 8723 6752
rect 8665 6743 8723 6749
rect 9030 6740 9036 6752
rect 9088 6740 9094 6792
rect 8021 6715 8079 6721
rect 8021 6712 8033 6715
rect 5552 6684 7328 6712
rect 7668 6684 8033 6712
rect 7668 6656 7696 6684
rect 8021 6681 8033 6684
rect 8067 6712 8079 6715
rect 8110 6712 8116 6724
rect 8067 6684 8116 6712
rect 8067 6681 8079 6684
rect 8021 6675 8079 6681
rect 8110 6672 8116 6684
rect 8168 6672 8174 6724
rect 4120 6616 5120 6644
rect 4120 6604 4126 6616
rect 5166 6604 5172 6656
rect 5224 6644 5230 6656
rect 5442 6644 5448 6656
rect 5224 6616 5448 6644
rect 5224 6604 5230 6616
rect 5442 6604 5448 6616
rect 5500 6644 5506 6656
rect 6454 6644 6460 6656
rect 5500 6616 6460 6644
rect 5500 6604 5506 6616
rect 6454 6604 6460 6616
rect 6512 6604 6518 6656
rect 7006 6604 7012 6656
rect 7064 6644 7070 6656
rect 7285 6647 7343 6653
rect 7285 6644 7297 6647
rect 7064 6616 7297 6644
rect 7064 6604 7070 6616
rect 7285 6613 7297 6616
rect 7331 6613 7343 6647
rect 7285 6607 7343 6613
rect 7466 6604 7472 6656
rect 7524 6604 7530 6656
rect 7650 6604 7656 6656
rect 7708 6604 7714 6656
rect 7742 6604 7748 6656
rect 7800 6644 7806 6656
rect 7837 6647 7895 6653
rect 7837 6644 7849 6647
rect 7800 6616 7849 6644
rect 7800 6604 7806 6616
rect 7837 6613 7849 6616
rect 7883 6613 7895 6647
rect 7837 6607 7895 6613
rect 8386 6604 8392 6656
rect 8444 6644 8450 6656
rect 8481 6647 8539 6653
rect 8481 6644 8493 6647
rect 8444 6616 8493 6644
rect 8444 6604 8450 6616
rect 8481 6613 8493 6616
rect 8527 6613 8539 6647
rect 8481 6607 8539 6613
rect 1104 6554 9016 6576
rect 1104 6502 2599 6554
rect 2651 6502 2663 6554
rect 2715 6502 2727 6554
rect 2779 6502 2791 6554
rect 2843 6502 2855 6554
rect 2907 6502 4577 6554
rect 4629 6502 4641 6554
rect 4693 6502 4705 6554
rect 4757 6502 4769 6554
rect 4821 6502 4833 6554
rect 4885 6502 6555 6554
rect 6607 6502 6619 6554
rect 6671 6502 6683 6554
rect 6735 6502 6747 6554
rect 6799 6502 6811 6554
rect 6863 6502 8533 6554
rect 8585 6502 8597 6554
rect 8649 6502 8661 6554
rect 8713 6502 8725 6554
rect 8777 6502 8789 6554
rect 8841 6502 9016 6554
rect 1104 6480 9016 6502
rect 2406 6440 2412 6452
rect 2240 6412 2412 6440
rect 1394 6332 1400 6384
rect 1452 6372 1458 6384
rect 2240 6381 2268 6412
rect 2406 6400 2412 6412
rect 2464 6400 2470 6452
rect 2498 6400 2504 6452
rect 2556 6400 2562 6452
rect 3326 6440 3332 6452
rect 2700 6412 3332 6440
rect 2700 6381 2728 6412
rect 3326 6400 3332 6412
rect 3384 6400 3390 6452
rect 4706 6440 4712 6452
rect 4172 6412 4712 6440
rect 2133 6375 2191 6381
rect 2133 6372 2145 6375
rect 1452 6344 2145 6372
rect 1452 6332 1458 6344
rect 2133 6341 2145 6344
rect 2179 6341 2191 6375
rect 2133 6335 2191 6341
rect 2225 6375 2283 6381
rect 2225 6341 2237 6375
rect 2271 6341 2283 6375
rect 2225 6335 2283 6341
rect 2685 6375 2743 6381
rect 2685 6341 2697 6375
rect 2731 6341 2743 6375
rect 2958 6372 2964 6384
rect 2685 6335 2743 6341
rect 2792 6344 2964 6372
rect 1581 6307 1639 6313
rect 1581 6273 1593 6307
rect 1627 6304 1639 6307
rect 1762 6304 1768 6316
rect 1627 6276 1768 6304
rect 1627 6273 1639 6276
rect 1581 6267 1639 6273
rect 1762 6264 1768 6276
rect 1820 6264 1826 6316
rect 1949 6307 2007 6313
rect 1949 6273 1961 6307
rect 1995 6304 2007 6307
rect 1995 6276 2268 6304
rect 1995 6273 2007 6276
rect 1949 6267 2007 6273
rect 1857 6239 1915 6245
rect 1857 6205 1869 6239
rect 1903 6236 1915 6239
rect 2240 6236 2268 6276
rect 2314 6264 2320 6316
rect 2372 6264 2378 6316
rect 2792 6236 2820 6344
rect 2958 6332 2964 6344
rect 3016 6332 3022 6384
rect 3602 6332 3608 6384
rect 3660 6372 3666 6384
rect 3660 6344 4108 6372
rect 3660 6332 3666 6344
rect 3050 6264 3056 6316
rect 3108 6304 3114 6316
rect 3237 6307 3295 6313
rect 3237 6304 3249 6307
rect 3108 6276 3249 6304
rect 3108 6264 3114 6276
rect 3237 6273 3249 6276
rect 3283 6273 3295 6307
rect 3237 6267 3295 6273
rect 3510 6264 3516 6316
rect 3568 6264 3574 6316
rect 3789 6307 3847 6313
rect 3789 6273 3801 6307
rect 3835 6304 3847 6307
rect 3878 6304 3884 6316
rect 3835 6276 3884 6304
rect 3835 6273 3847 6276
rect 3789 6267 3847 6273
rect 3878 6264 3884 6276
rect 3936 6264 3942 6316
rect 3970 6264 3976 6316
rect 4028 6264 4034 6316
rect 1903 6208 2176 6236
rect 2240 6208 2820 6236
rect 3145 6239 3203 6245
rect 1903 6205 1915 6208
rect 1857 6199 1915 6205
rect 1394 6060 1400 6112
rect 1452 6060 1458 6112
rect 1762 6060 1768 6112
rect 1820 6060 1826 6112
rect 2148 6100 2176 6208
rect 3145 6205 3157 6239
rect 3191 6236 3203 6239
rect 3988 6236 4016 6264
rect 3191 6208 4016 6236
rect 4080 6236 4108 6344
rect 4172 6313 4200 6412
rect 4706 6400 4712 6412
rect 4764 6440 4770 6452
rect 7101 6443 7159 6449
rect 4764 6412 5856 6440
rect 4764 6400 4770 6412
rect 5828 6384 5856 6412
rect 7101 6409 7113 6443
rect 7147 6440 7159 6443
rect 7374 6440 7380 6452
rect 7147 6412 7380 6440
rect 7147 6409 7159 6412
rect 7101 6403 7159 6409
rect 7374 6400 7380 6412
rect 7432 6400 7438 6452
rect 7466 6400 7472 6452
rect 7524 6400 7530 6452
rect 4433 6375 4491 6381
rect 4433 6372 4445 6375
rect 4264 6344 4445 6372
rect 4157 6307 4215 6313
rect 4157 6273 4169 6307
rect 4203 6273 4215 6307
rect 4157 6267 4215 6273
rect 4264 6236 4292 6344
rect 4433 6341 4445 6344
rect 4479 6341 4491 6375
rect 4433 6335 4491 6341
rect 5626 6332 5632 6384
rect 5684 6332 5690 6384
rect 5810 6332 5816 6384
rect 5868 6332 5874 6384
rect 6178 6332 6184 6384
rect 6236 6372 6242 6384
rect 6236 6344 6684 6372
rect 6236 6332 6242 6344
rect 4341 6307 4399 6313
rect 4341 6273 4353 6307
rect 4387 6304 4399 6307
rect 4522 6304 4528 6316
rect 4387 6276 4528 6304
rect 4387 6273 4399 6276
rect 4341 6267 4399 6273
rect 4522 6264 4528 6276
rect 4580 6304 4586 6316
rect 5644 6304 5672 6332
rect 4580 6276 5672 6304
rect 4580 6264 4586 6276
rect 5718 6264 5724 6316
rect 5776 6304 5782 6316
rect 6362 6304 6368 6316
rect 5776 6276 6368 6304
rect 5776 6264 5782 6276
rect 6362 6264 6368 6276
rect 6420 6264 6426 6316
rect 6656 6313 6684 6344
rect 6641 6307 6699 6313
rect 6641 6273 6653 6307
rect 6687 6273 6699 6307
rect 6641 6267 6699 6273
rect 6914 6264 6920 6316
rect 6972 6264 6978 6316
rect 7282 6264 7288 6316
rect 7340 6264 7346 6316
rect 7484 6304 7512 6400
rect 7541 6307 7599 6313
rect 7541 6304 7553 6307
rect 7484 6276 7553 6304
rect 7541 6273 7553 6276
rect 7587 6273 7599 6307
rect 7541 6267 7599 6273
rect 4080 6208 4292 6236
rect 7193 6239 7251 6245
rect 3191 6205 3203 6208
rect 3145 6199 3203 6205
rect 7193 6205 7205 6239
rect 7239 6205 7251 6239
rect 7193 6199 7251 6205
rect 2222 6128 2228 6180
rect 2280 6168 2286 6180
rect 2961 6171 3019 6177
rect 2961 6168 2973 6171
rect 2280 6140 2973 6168
rect 2280 6128 2286 6140
rect 2961 6137 2973 6140
rect 3007 6137 3019 6171
rect 2961 6131 3019 6137
rect 3326 6100 3332 6112
rect 2148 6072 3332 6100
rect 3326 6060 3332 6072
rect 3384 6060 3390 6112
rect 3602 6060 3608 6112
rect 3660 6100 3666 6112
rect 4062 6100 4068 6112
rect 3660 6072 4068 6100
rect 3660 6060 3666 6072
rect 4062 6060 4068 6072
rect 4120 6060 4126 6112
rect 4338 6060 4344 6112
rect 4396 6100 4402 6112
rect 5721 6103 5779 6109
rect 5721 6100 5733 6103
rect 4396 6072 5733 6100
rect 4396 6060 4402 6072
rect 5721 6069 5733 6072
rect 5767 6069 5779 6103
rect 5721 6063 5779 6069
rect 6454 6060 6460 6112
rect 6512 6100 6518 6112
rect 7208 6100 7236 6199
rect 7282 6100 7288 6112
rect 6512 6072 7288 6100
rect 6512 6060 6518 6072
rect 7282 6060 7288 6072
rect 7340 6100 7346 6112
rect 7926 6100 7932 6112
rect 7340 6072 7932 6100
rect 7340 6060 7346 6072
rect 7926 6060 7932 6072
rect 7984 6060 7990 6112
rect 8665 6103 8723 6109
rect 8665 6069 8677 6103
rect 8711 6100 8723 6103
rect 8938 6100 8944 6112
rect 8711 6072 8944 6100
rect 8711 6069 8723 6072
rect 8665 6063 8723 6069
rect 8938 6060 8944 6072
rect 8996 6060 9002 6112
rect 1104 6010 9016 6032
rect 1104 5958 1939 6010
rect 1991 5958 2003 6010
rect 2055 5958 2067 6010
rect 2119 5958 2131 6010
rect 2183 5958 2195 6010
rect 2247 5958 3917 6010
rect 3969 5958 3981 6010
rect 4033 5958 4045 6010
rect 4097 5958 4109 6010
rect 4161 5958 4173 6010
rect 4225 5958 5895 6010
rect 5947 5958 5959 6010
rect 6011 5958 6023 6010
rect 6075 5958 6087 6010
rect 6139 5958 6151 6010
rect 6203 5958 7873 6010
rect 7925 5958 7937 6010
rect 7989 5958 8001 6010
rect 8053 5958 8065 6010
rect 8117 5958 8129 6010
rect 8181 5958 9016 6010
rect 1104 5936 9016 5958
rect 1394 5856 1400 5908
rect 1452 5856 1458 5908
rect 1581 5899 1639 5905
rect 1581 5865 1593 5899
rect 1627 5896 1639 5899
rect 1670 5896 1676 5908
rect 1627 5868 1676 5896
rect 1627 5865 1639 5868
rect 1581 5859 1639 5865
rect 1670 5856 1676 5868
rect 1728 5856 1734 5908
rect 1762 5856 1768 5908
rect 1820 5896 1826 5908
rect 2225 5899 2283 5905
rect 2225 5896 2237 5899
rect 1820 5868 2237 5896
rect 1820 5856 1826 5868
rect 2225 5865 2237 5868
rect 2271 5865 2283 5899
rect 4614 5896 4620 5908
rect 2225 5859 2283 5865
rect 3712 5868 4620 5896
rect 1412 5692 1440 5856
rect 3712 5828 3740 5868
rect 4614 5856 4620 5868
rect 4672 5856 4678 5908
rect 4985 5899 5043 5905
rect 4985 5865 4997 5899
rect 5031 5865 5043 5899
rect 5534 5896 5540 5908
rect 4985 5859 5043 5865
rect 5368 5868 5540 5896
rect 2240 5800 3740 5828
rect 3789 5831 3847 5837
rect 2240 5704 2268 5800
rect 3789 5797 3801 5831
rect 3835 5828 3847 5831
rect 5000 5828 5028 5859
rect 5368 5828 5396 5868
rect 5534 5856 5540 5868
rect 5592 5856 5598 5908
rect 5994 5856 6000 5908
rect 6052 5896 6058 5908
rect 6089 5899 6147 5905
rect 6089 5896 6101 5899
rect 6052 5868 6101 5896
rect 6052 5856 6058 5868
rect 6089 5865 6101 5868
rect 6135 5865 6147 5899
rect 6089 5859 6147 5865
rect 7006 5856 7012 5908
rect 7064 5856 7070 5908
rect 7558 5856 7564 5908
rect 7616 5856 7622 5908
rect 7742 5856 7748 5908
rect 7800 5856 7806 5908
rect 8021 5899 8079 5905
rect 8021 5865 8033 5899
rect 8067 5896 8079 5899
rect 8202 5896 8208 5908
rect 8067 5868 8208 5896
rect 8067 5865 8079 5868
rect 8021 5859 8079 5865
rect 8202 5856 8208 5868
rect 8260 5856 8266 5908
rect 5810 5828 5816 5840
rect 3835 5800 4200 5828
rect 5000 5800 5396 5828
rect 3835 5797 3847 5800
rect 3789 5791 3847 5797
rect 3329 5763 3387 5769
rect 3329 5760 3341 5763
rect 2332 5732 3341 5760
rect 2332 5704 2360 5732
rect 3329 5729 3341 5732
rect 3375 5760 3387 5763
rect 3694 5760 3700 5772
rect 3375 5732 3700 5760
rect 3375 5729 3387 5732
rect 3329 5723 3387 5729
rect 3694 5720 3700 5732
rect 3752 5720 3758 5772
rect 4172 5704 4200 5800
rect 4798 5760 4804 5772
rect 4632 5732 4804 5760
rect 1765 5695 1823 5701
rect 1765 5692 1777 5695
rect 1412 5664 1777 5692
rect 1765 5661 1777 5664
rect 1811 5661 1823 5695
rect 1765 5655 1823 5661
rect 1854 5652 1860 5704
rect 1912 5692 1918 5704
rect 1949 5695 2007 5701
rect 1949 5692 1961 5695
rect 1912 5664 1961 5692
rect 1912 5652 1918 5664
rect 1949 5661 1961 5664
rect 1995 5661 2007 5695
rect 1949 5655 2007 5661
rect 2041 5695 2099 5701
rect 2041 5661 2053 5695
rect 2087 5692 2099 5695
rect 2222 5692 2228 5704
rect 2087 5664 2228 5692
rect 2087 5661 2099 5664
rect 2041 5655 2099 5661
rect 2222 5652 2228 5664
rect 2280 5652 2286 5704
rect 2314 5652 2320 5704
rect 2372 5652 2378 5704
rect 2409 5695 2467 5701
rect 2409 5661 2421 5695
rect 2455 5661 2467 5695
rect 2409 5655 2467 5661
rect 2424 5624 2452 5655
rect 2498 5652 2504 5704
rect 2556 5692 2562 5704
rect 2593 5695 2651 5701
rect 2593 5692 2605 5695
rect 2556 5664 2605 5692
rect 2556 5652 2562 5664
rect 2593 5661 2605 5664
rect 2639 5661 2651 5695
rect 2593 5655 2651 5661
rect 2685 5695 2743 5701
rect 2685 5661 2697 5695
rect 2731 5692 2743 5695
rect 2866 5692 2872 5704
rect 2731 5664 2872 5692
rect 2731 5661 2743 5664
rect 2685 5655 2743 5661
rect 2866 5652 2872 5664
rect 2924 5652 2930 5704
rect 3510 5692 3516 5704
rect 2971 5664 3516 5692
rect 2971 5624 2999 5664
rect 3510 5652 3516 5664
rect 3568 5652 3574 5704
rect 3620 5664 3924 5692
rect 2424 5596 2999 5624
rect 3234 5584 3240 5636
rect 3292 5624 3298 5636
rect 3620 5624 3648 5664
rect 3896 5633 3924 5664
rect 3970 5652 3976 5704
rect 4028 5652 4034 5704
rect 4062 5652 4068 5704
rect 4120 5652 4126 5704
rect 4154 5652 4160 5704
rect 4212 5652 4218 5704
rect 4246 5652 4252 5704
rect 4304 5652 4310 5704
rect 4632 5701 4660 5732
rect 4798 5720 4804 5732
rect 4856 5720 4862 5772
rect 5077 5763 5135 5769
rect 5077 5729 5089 5763
rect 5123 5729 5135 5763
rect 5077 5726 5135 5729
rect 5031 5723 5135 5726
rect 5031 5704 5120 5723
rect 4617 5695 4675 5701
rect 4617 5661 4629 5695
rect 4663 5661 4675 5695
rect 4617 5655 4675 5661
rect 4706 5652 4712 5704
rect 4764 5692 4770 5704
rect 4893 5695 4951 5701
rect 4893 5692 4905 5695
rect 4764 5664 4905 5692
rect 4764 5652 4770 5664
rect 4893 5661 4905 5664
rect 4939 5661 4951 5695
rect 4893 5655 4951 5661
rect 4982 5652 4988 5704
rect 5040 5698 5120 5704
rect 5040 5652 5059 5698
rect 5166 5652 5172 5704
rect 5224 5652 5230 5704
rect 5368 5692 5396 5800
rect 5552 5800 5816 5828
rect 5442 5720 5448 5772
rect 5500 5760 5506 5772
rect 5552 5769 5580 5800
rect 5810 5788 5816 5800
rect 5868 5788 5874 5840
rect 6454 5828 6460 5840
rect 6380 5800 6460 5828
rect 5537 5763 5595 5769
rect 5537 5760 5549 5763
rect 5500 5732 5549 5760
rect 5500 5720 5506 5732
rect 5537 5729 5549 5732
rect 5583 5729 5595 5763
rect 5537 5723 5595 5729
rect 5626 5720 5632 5772
rect 5684 5760 5690 5772
rect 5721 5763 5779 5769
rect 5721 5760 5733 5763
rect 5684 5732 5733 5760
rect 5684 5720 5690 5732
rect 5721 5729 5733 5732
rect 5767 5760 5779 5763
rect 6380 5760 6408 5800
rect 6454 5788 6460 5800
rect 6512 5788 6518 5840
rect 6917 5831 6975 5837
rect 6917 5797 6929 5831
rect 6963 5828 6975 5831
rect 7576 5828 7604 5856
rect 6963 5800 7604 5828
rect 6963 5797 6975 5800
rect 6917 5791 6975 5797
rect 7760 5769 7788 5856
rect 8386 5828 8392 5840
rect 8220 5800 8392 5828
rect 6733 5763 6791 5769
rect 6733 5760 6745 5763
rect 5767 5732 6408 5760
rect 5767 5729 5779 5732
rect 5721 5723 5779 5729
rect 6380 5701 6408 5732
rect 6472 5732 6745 5760
rect 6472 5704 6500 5732
rect 6733 5729 6745 5732
rect 6779 5729 6791 5763
rect 6733 5723 6791 5729
rect 7745 5763 7803 5769
rect 7745 5729 7757 5763
rect 7791 5729 7803 5763
rect 7745 5723 7803 5729
rect 8220 5704 8248 5800
rect 8386 5788 8392 5800
rect 8444 5788 8450 5840
rect 5813 5695 5871 5701
rect 5813 5692 5825 5695
rect 5368 5664 5825 5692
rect 5813 5661 5825 5664
rect 5859 5661 5871 5695
rect 5813 5655 5871 5661
rect 6365 5695 6423 5701
rect 6365 5661 6377 5695
rect 6411 5661 6423 5695
rect 6365 5655 6423 5661
rect 3292 5596 3648 5624
rect 3881 5627 3939 5633
rect 3292 5584 3298 5596
rect 3881 5593 3893 5627
rect 3927 5593 3939 5627
rect 3988 5624 4016 5652
rect 5031 5624 5059 5652
rect 3988 5596 5059 5624
rect 5828 5624 5856 5655
rect 6454 5652 6460 5704
rect 6512 5652 6518 5704
rect 6549 5695 6607 5701
rect 6549 5661 6561 5695
rect 6595 5661 6607 5695
rect 6549 5655 6607 5661
rect 6564 5624 6592 5655
rect 6914 5652 6920 5704
rect 6972 5652 6978 5704
rect 7006 5652 7012 5704
rect 7064 5692 7070 5704
rect 7190 5692 7196 5704
rect 7064 5664 7196 5692
rect 7064 5652 7070 5664
rect 7190 5652 7196 5664
rect 7248 5692 7254 5704
rect 7285 5695 7343 5701
rect 7285 5692 7297 5695
rect 7248 5664 7297 5692
rect 7248 5652 7254 5664
rect 7285 5661 7297 5664
rect 7331 5661 7343 5695
rect 7285 5655 7343 5661
rect 7650 5652 7656 5704
rect 7708 5652 7714 5704
rect 8202 5652 8208 5704
rect 8260 5652 8266 5704
rect 8386 5652 8392 5704
rect 8444 5692 8450 5704
rect 8573 5695 8631 5701
rect 8573 5692 8585 5695
rect 8444 5664 8585 5692
rect 8444 5652 8450 5664
rect 8573 5661 8585 5664
rect 8619 5661 8631 5695
rect 8573 5655 8631 5661
rect 5828 5596 7512 5624
rect 3881 5587 3939 5593
rect 7484 5568 7512 5596
rect 1578 5516 1584 5568
rect 1636 5556 1642 5568
rect 2498 5556 2504 5568
rect 1636 5528 2504 5556
rect 1636 5516 1642 5528
rect 2498 5516 2504 5528
rect 2556 5516 2562 5568
rect 2777 5559 2835 5565
rect 2777 5525 2789 5559
rect 2823 5556 2835 5559
rect 2958 5556 2964 5568
rect 2823 5528 2964 5556
rect 2823 5525 2835 5528
rect 2777 5519 2835 5525
rect 2958 5516 2964 5528
rect 3016 5516 3022 5568
rect 4154 5516 4160 5568
rect 4212 5556 4218 5568
rect 4709 5559 4767 5565
rect 4709 5556 4721 5559
rect 4212 5528 4721 5556
rect 4212 5516 4218 5528
rect 4709 5525 4721 5528
rect 4755 5525 4767 5559
rect 4709 5519 4767 5525
rect 4798 5516 4804 5568
rect 4856 5556 4862 5568
rect 5350 5556 5356 5568
rect 4856 5528 5356 5556
rect 4856 5516 4862 5528
rect 5350 5516 5356 5528
rect 5408 5516 5414 5568
rect 5626 5516 5632 5568
rect 5684 5556 5690 5568
rect 5905 5559 5963 5565
rect 5905 5556 5917 5559
rect 5684 5528 5917 5556
rect 5684 5516 5690 5528
rect 5905 5525 5917 5528
rect 5951 5525 5963 5559
rect 5905 5519 5963 5525
rect 6270 5516 6276 5568
rect 6328 5556 6334 5568
rect 6641 5559 6699 5565
rect 6641 5556 6653 5559
rect 6328 5528 6653 5556
rect 6328 5516 6334 5528
rect 6641 5525 6653 5528
rect 6687 5556 6699 5559
rect 7377 5559 7435 5565
rect 7377 5556 7389 5559
rect 6687 5528 7389 5556
rect 6687 5525 6699 5528
rect 6641 5519 6699 5525
rect 7377 5525 7389 5528
rect 7423 5525 7435 5559
rect 7377 5519 7435 5525
rect 7466 5516 7472 5568
rect 7524 5516 7530 5568
rect 1104 5466 9016 5488
rect 1104 5414 2599 5466
rect 2651 5414 2663 5466
rect 2715 5414 2727 5466
rect 2779 5414 2791 5466
rect 2843 5414 2855 5466
rect 2907 5414 4577 5466
rect 4629 5414 4641 5466
rect 4693 5414 4705 5466
rect 4757 5414 4769 5466
rect 4821 5414 4833 5466
rect 4885 5414 6555 5466
rect 6607 5414 6619 5466
rect 6671 5414 6683 5466
rect 6735 5414 6747 5466
rect 6799 5414 6811 5466
rect 6863 5414 8533 5466
rect 8585 5414 8597 5466
rect 8649 5414 8661 5466
rect 8713 5414 8725 5466
rect 8777 5414 8789 5466
rect 8841 5414 9016 5466
rect 1104 5392 9016 5414
rect 2866 5312 2872 5364
rect 2924 5352 2930 5364
rect 3145 5355 3203 5361
rect 3145 5352 3157 5355
rect 2924 5324 3157 5352
rect 2924 5312 2930 5324
rect 3145 5321 3157 5324
rect 3191 5352 3203 5355
rect 3697 5355 3755 5361
rect 3697 5352 3709 5355
rect 3191 5324 3709 5352
rect 3191 5321 3203 5324
rect 3145 5315 3203 5321
rect 3697 5321 3709 5324
rect 3743 5321 3755 5355
rect 3697 5315 3755 5321
rect 4062 5312 4068 5364
rect 4120 5352 4126 5364
rect 4614 5352 4620 5364
rect 4120 5324 4620 5352
rect 4120 5312 4126 5324
rect 3050 5244 3056 5296
rect 3108 5244 3114 5296
rect 3234 5244 3240 5296
rect 3292 5244 3298 5296
rect 1664 5219 1722 5225
rect 1664 5185 1676 5219
rect 1710 5216 1722 5219
rect 2869 5219 2927 5225
rect 1710 5188 2452 5216
rect 1710 5185 1722 5188
rect 1664 5179 1722 5185
rect 1394 5108 1400 5160
rect 1452 5108 1458 5160
rect 2424 5080 2452 5188
rect 2869 5185 2881 5219
rect 2915 5216 2927 5219
rect 2958 5216 2964 5228
rect 2915 5188 2964 5216
rect 2915 5185 2927 5188
rect 2869 5179 2927 5185
rect 2958 5176 2964 5188
rect 3016 5176 3022 5228
rect 3068 5157 3096 5244
rect 3329 5219 3387 5225
rect 3329 5185 3341 5219
rect 3375 5185 3387 5219
rect 3329 5179 3387 5185
rect 3053 5151 3111 5157
rect 3053 5117 3065 5151
rect 3099 5117 3111 5151
rect 3053 5111 3111 5117
rect 2961 5083 3019 5089
rect 2961 5080 2973 5083
rect 2424 5052 2973 5080
rect 2961 5049 2973 5052
rect 3007 5049 3019 5083
rect 3344 5080 3372 5179
rect 3694 5176 3700 5228
rect 3752 5216 3758 5228
rect 4172 5216 4200 5324
rect 4614 5312 4620 5324
rect 4672 5312 4678 5364
rect 4706 5312 4712 5364
rect 4764 5352 4770 5364
rect 4764 5324 4844 5352
rect 4764 5312 4770 5324
rect 4246 5244 4252 5296
rect 4304 5284 4310 5296
rect 4816 5284 4844 5324
rect 5350 5312 5356 5364
rect 5408 5352 5414 5364
rect 6362 5352 6368 5364
rect 5408 5324 6368 5352
rect 5408 5312 5414 5324
rect 6362 5312 6368 5324
rect 6420 5352 6426 5364
rect 6825 5355 6883 5361
rect 6825 5352 6837 5355
rect 6420 5324 6837 5352
rect 6420 5312 6426 5324
rect 6825 5321 6837 5324
rect 6871 5321 6883 5355
rect 6825 5315 6883 5321
rect 6914 5312 6920 5364
rect 6972 5312 6978 5364
rect 7377 5355 7435 5361
rect 7377 5321 7389 5355
rect 7423 5352 7435 5355
rect 7466 5352 7472 5364
rect 7423 5324 7472 5352
rect 7423 5321 7435 5324
rect 7377 5315 7435 5321
rect 7466 5312 7472 5324
rect 7524 5312 7530 5364
rect 8573 5355 8631 5361
rect 8573 5352 8585 5355
rect 8036 5324 8585 5352
rect 5442 5284 5448 5296
rect 4304 5256 4752 5284
rect 4816 5256 5448 5284
rect 4304 5244 4310 5256
rect 3752 5188 4200 5216
rect 3752 5176 3758 5188
rect 4430 5176 4436 5228
rect 4488 5216 4494 5228
rect 4724 5225 4752 5256
rect 5442 5244 5448 5256
rect 5500 5244 5506 5296
rect 5718 5244 5724 5296
rect 5776 5284 5782 5296
rect 6932 5284 6960 5312
rect 7558 5284 7564 5296
rect 5776 5256 6040 5284
rect 6932 5256 7564 5284
rect 5776 5244 5782 5256
rect 4709 5219 4767 5225
rect 4488 5188 4660 5216
rect 4488 5176 4494 5188
rect 3513 5151 3571 5157
rect 3513 5117 3525 5151
rect 3559 5148 3571 5151
rect 3878 5148 3884 5160
rect 3559 5120 3884 5148
rect 3559 5117 3571 5120
rect 3513 5111 3571 5117
rect 3878 5108 3884 5120
rect 3936 5108 3942 5160
rect 4065 5151 4123 5157
rect 4065 5117 4077 5151
rect 4111 5148 4123 5151
rect 4246 5148 4252 5160
rect 4111 5120 4252 5148
rect 4111 5117 4123 5120
rect 4065 5111 4123 5117
rect 4246 5108 4252 5120
rect 4304 5108 4310 5160
rect 4341 5151 4399 5157
rect 4341 5117 4353 5151
rect 4387 5148 4399 5151
rect 4632 5148 4660 5188
rect 4709 5185 4721 5219
rect 4755 5216 4767 5219
rect 4798 5216 4804 5228
rect 4755 5188 4804 5216
rect 4755 5185 4767 5188
rect 4709 5179 4767 5185
rect 4798 5176 4804 5188
rect 4856 5176 4862 5228
rect 5077 5219 5135 5225
rect 5077 5185 5089 5219
rect 5123 5216 5135 5219
rect 5350 5216 5356 5228
rect 5123 5188 5356 5216
rect 5123 5185 5135 5188
rect 5077 5179 5135 5185
rect 5350 5176 5356 5188
rect 5408 5176 5414 5228
rect 5460 5216 5488 5244
rect 5537 5219 5595 5225
rect 5537 5216 5549 5219
rect 5460 5188 5549 5216
rect 5537 5185 5549 5188
rect 5583 5185 5595 5219
rect 5537 5179 5595 5185
rect 5626 5176 5632 5228
rect 5684 5176 5690 5228
rect 6012 5225 6040 5256
rect 7558 5244 7564 5256
rect 7616 5284 7622 5296
rect 8036 5284 8064 5324
rect 8573 5321 8585 5324
rect 8619 5321 8631 5355
rect 8573 5315 8631 5321
rect 7616 5256 8064 5284
rect 7616 5244 7622 5256
rect 8294 5244 8300 5296
rect 8352 5284 8358 5296
rect 8352 5256 8708 5284
rect 8352 5244 8358 5256
rect 5813 5219 5871 5225
rect 5813 5185 5825 5219
rect 5859 5185 5871 5219
rect 5813 5179 5871 5185
rect 5997 5219 6055 5225
rect 5997 5185 6009 5219
rect 6043 5185 6055 5219
rect 5997 5179 6055 5185
rect 5721 5151 5779 5157
rect 5721 5148 5733 5151
rect 4387 5120 4568 5148
rect 4632 5120 5733 5148
rect 4387 5117 4399 5120
rect 4341 5111 4399 5117
rect 4154 5080 4160 5092
rect 3344 5052 4160 5080
rect 2961 5043 3019 5049
rect 4154 5040 4160 5052
rect 4212 5040 4218 5092
rect 1762 4972 1768 5024
rect 1820 5012 1826 5024
rect 2590 5012 2596 5024
rect 1820 4984 2596 5012
rect 1820 4972 1826 4984
rect 2590 4972 2596 4984
rect 2648 4972 2654 5024
rect 2777 5015 2835 5021
rect 2777 4981 2789 5015
rect 2823 5012 2835 5015
rect 3970 5012 3976 5024
rect 2823 4984 3976 5012
rect 2823 4981 2835 4984
rect 2777 4975 2835 4981
rect 3970 4972 3976 4984
rect 4028 4972 4034 5024
rect 4540 5012 4568 5120
rect 5721 5117 5733 5120
rect 5767 5117 5779 5151
rect 5828 5148 5856 5179
rect 6178 5176 6184 5228
rect 6236 5176 6242 5228
rect 6638 5176 6644 5228
rect 6696 5216 6702 5228
rect 7101 5219 7159 5225
rect 7101 5216 7113 5219
rect 6696 5188 7113 5216
rect 6696 5176 6702 5188
rect 7101 5185 7113 5188
rect 7147 5185 7159 5219
rect 8202 5216 8208 5228
rect 7101 5179 7159 5185
rect 7556 5188 8208 5216
rect 6196 5148 6224 5176
rect 5828 5120 6224 5148
rect 6365 5151 6423 5157
rect 5721 5111 5779 5117
rect 6365 5117 6377 5151
rect 6411 5148 6423 5151
rect 7556 5148 7584 5188
rect 8202 5176 8208 5188
rect 8260 5176 8266 5228
rect 8386 5176 8392 5228
rect 8444 5176 8450 5228
rect 8680 5225 8708 5256
rect 8665 5219 8723 5225
rect 8665 5185 8677 5219
rect 8711 5185 8723 5219
rect 8665 5179 8723 5185
rect 6411 5120 7584 5148
rect 6411 5117 6423 5120
rect 6365 5111 6423 5117
rect 4982 5040 4988 5092
rect 5040 5040 5046 5092
rect 5074 5040 5080 5092
rect 5132 5080 5138 5092
rect 5810 5080 5816 5092
rect 5132 5052 5816 5080
rect 5132 5040 5138 5052
rect 5810 5040 5816 5052
rect 5868 5040 5874 5092
rect 6380 5080 6408 5111
rect 7650 5108 7656 5160
rect 7708 5108 7714 5160
rect 7742 5108 7748 5160
rect 7800 5148 7806 5160
rect 8113 5151 8171 5157
rect 8113 5148 8125 5151
rect 7800 5120 8125 5148
rect 7800 5108 7806 5120
rect 8113 5117 8125 5120
rect 8159 5117 8171 5151
rect 8113 5111 8171 5117
rect 5920 5052 6408 5080
rect 5092 5012 5120 5040
rect 4540 4984 5120 5012
rect 5350 4972 5356 5024
rect 5408 4972 5414 5024
rect 5442 4972 5448 5024
rect 5500 5012 5506 5024
rect 5920 5012 5948 5052
rect 6638 5040 6644 5092
rect 6696 5040 6702 5092
rect 7668 5080 7696 5108
rect 8389 5083 8447 5089
rect 8389 5080 8401 5083
rect 7668 5052 8401 5080
rect 8389 5049 8401 5052
rect 8435 5049 8447 5083
rect 8389 5043 8447 5049
rect 5500 4984 5948 5012
rect 5500 4972 5506 4984
rect 5994 4972 6000 5024
rect 6052 5012 6058 5024
rect 6730 5012 6736 5024
rect 6052 4984 6736 5012
rect 6052 4972 6058 4984
rect 6730 4972 6736 4984
rect 6788 4972 6794 5024
rect 7558 4972 7564 5024
rect 7616 4972 7622 5024
rect 1104 4922 9016 4944
rect 1104 4870 1939 4922
rect 1991 4870 2003 4922
rect 2055 4870 2067 4922
rect 2119 4870 2131 4922
rect 2183 4870 2195 4922
rect 2247 4870 3917 4922
rect 3969 4870 3981 4922
rect 4033 4870 4045 4922
rect 4097 4870 4109 4922
rect 4161 4870 4173 4922
rect 4225 4870 5895 4922
rect 5947 4870 5959 4922
rect 6011 4870 6023 4922
rect 6075 4870 6087 4922
rect 6139 4870 6151 4922
rect 6203 4870 7873 4922
rect 7925 4870 7937 4922
rect 7989 4870 8001 4922
rect 8053 4870 8065 4922
rect 8117 4870 8129 4922
rect 8181 4870 9016 4922
rect 1104 4848 9016 4870
rect 1762 4768 1768 4820
rect 1820 4768 1826 4820
rect 1857 4811 1915 4817
rect 1857 4777 1869 4811
rect 1903 4808 1915 4811
rect 3050 4808 3056 4820
rect 1903 4780 3056 4808
rect 1903 4777 1915 4780
rect 1857 4771 1915 4777
rect 3050 4768 3056 4780
rect 3108 4768 3114 4820
rect 3142 4768 3148 4820
rect 3200 4808 3206 4820
rect 3200 4780 3648 4808
rect 3200 4768 3206 4780
rect 1581 4607 1639 4613
rect 1581 4573 1593 4607
rect 1627 4604 1639 4607
rect 1780 4604 1808 4768
rect 3421 4743 3479 4749
rect 2516 4712 3280 4740
rect 2314 4632 2320 4684
rect 2372 4632 2378 4684
rect 2516 4681 2544 4712
rect 3252 4681 3280 4712
rect 3421 4709 3433 4743
rect 3467 4740 3479 4743
rect 3510 4740 3516 4752
rect 3467 4712 3516 4740
rect 3467 4709 3479 4712
rect 3421 4703 3479 4709
rect 3510 4700 3516 4712
rect 3568 4700 3574 4752
rect 3620 4681 3648 4780
rect 3970 4768 3976 4820
rect 4028 4808 4034 4820
rect 5166 4808 5172 4820
rect 4028 4780 5172 4808
rect 4028 4768 4034 4780
rect 5166 4768 5172 4780
rect 5224 4768 5230 4820
rect 5368 4780 5764 4808
rect 5368 4740 5396 4780
rect 4356 4712 5396 4740
rect 4356 4681 4384 4712
rect 5442 4700 5448 4752
rect 5500 4740 5506 4752
rect 5736 4749 5764 4780
rect 6454 4768 6460 4820
rect 6512 4768 6518 4820
rect 6730 4768 6736 4820
rect 6788 4768 6794 4820
rect 7006 4768 7012 4820
rect 7064 4768 7070 4820
rect 7466 4768 7472 4820
rect 7524 4768 7530 4820
rect 8202 4768 8208 4820
rect 8260 4768 8266 4820
rect 5537 4743 5595 4749
rect 5537 4740 5549 4743
rect 5500 4712 5549 4740
rect 5500 4700 5506 4712
rect 5537 4709 5549 4712
rect 5583 4709 5595 4743
rect 5537 4703 5595 4709
rect 5721 4743 5779 4749
rect 5721 4709 5733 4743
rect 5767 4709 5779 4743
rect 7024 4740 7052 4768
rect 5721 4703 5779 4709
rect 6104 4712 7052 4740
rect 2501 4675 2559 4681
rect 2501 4641 2513 4675
rect 2547 4641 2559 4675
rect 2501 4635 2559 4641
rect 3237 4675 3295 4681
rect 3237 4641 3249 4675
rect 3283 4672 3295 4675
rect 3605 4675 3663 4681
rect 3283 4644 3464 4672
rect 3283 4641 3295 4644
rect 3237 4635 3295 4641
rect 3436 4616 3464 4644
rect 3605 4641 3617 4675
rect 3651 4641 3663 4675
rect 3605 4635 3663 4641
rect 4341 4675 4399 4681
rect 4341 4641 4353 4675
rect 4387 4641 4399 4675
rect 4341 4635 4399 4641
rect 4430 4632 4436 4684
rect 4488 4672 4494 4684
rect 4709 4675 4767 4681
rect 4488 4644 4660 4672
rect 4488 4632 4494 4644
rect 1627 4576 1808 4604
rect 1857 4607 1915 4613
rect 1627 4573 1639 4576
rect 1581 4567 1639 4573
rect 1857 4573 1869 4607
rect 1903 4604 1915 4607
rect 2041 4607 2099 4613
rect 2041 4604 2053 4607
rect 1903 4576 2053 4604
rect 1903 4573 1915 4576
rect 1857 4567 1915 4573
rect 2041 4573 2053 4576
rect 2087 4573 2099 4607
rect 2041 4567 2099 4573
rect 2225 4607 2283 4613
rect 2225 4573 2237 4607
rect 2271 4604 2283 4607
rect 3050 4604 3056 4616
rect 2271 4576 3056 4604
rect 2271 4573 2283 4576
rect 2225 4567 2283 4573
rect 1765 4539 1823 4545
rect 1765 4505 1777 4539
rect 1811 4505 1823 4539
rect 1765 4499 1823 4505
rect 1780 4468 1808 4499
rect 1946 4496 1952 4548
rect 2004 4496 2010 4548
rect 2056 4536 2084 4567
rect 3050 4564 3056 4576
rect 3108 4564 3114 4616
rect 3329 4607 3387 4613
rect 3329 4573 3341 4607
rect 3375 4573 3387 4607
rect 3329 4567 3387 4573
rect 2056 4508 2774 4536
rect 2130 4468 2136 4480
rect 1780 4440 2136 4468
rect 2130 4428 2136 4440
rect 2188 4428 2194 4480
rect 2590 4428 2596 4480
rect 2648 4428 2654 4480
rect 2746 4468 2774 4508
rect 2866 4496 2872 4548
rect 2924 4536 2930 4548
rect 3344 4536 3372 4567
rect 3418 4564 3424 4616
rect 3476 4564 3482 4616
rect 3973 4607 4031 4613
rect 3973 4573 3985 4607
rect 4019 4573 4031 4607
rect 3973 4567 4031 4573
rect 2924 4508 3372 4536
rect 3988 4536 4016 4567
rect 4062 4564 4068 4616
rect 4120 4564 4126 4616
rect 4157 4607 4215 4613
rect 4157 4573 4169 4607
rect 4203 4604 4215 4607
rect 4203 4576 4384 4604
rect 4203 4573 4215 4576
rect 4157 4567 4215 4573
rect 3988 4508 4108 4536
rect 2924 4496 2930 4508
rect 4080 4480 4108 4508
rect 3234 4468 3240 4480
rect 2746 4440 3240 4468
rect 3234 4428 3240 4440
rect 3292 4428 3298 4480
rect 3326 4428 3332 4480
rect 3384 4428 3390 4480
rect 4062 4428 4068 4480
rect 4120 4428 4126 4480
rect 4246 4428 4252 4480
rect 4304 4428 4310 4480
rect 4356 4468 4384 4576
rect 4522 4564 4528 4616
rect 4580 4564 4586 4616
rect 4632 4604 4660 4644
rect 4709 4641 4721 4675
rect 4755 4672 4767 4675
rect 5074 4672 5080 4684
rect 4755 4644 5080 4672
rect 4755 4641 4767 4644
rect 4709 4635 4767 4641
rect 5074 4632 5080 4644
rect 5132 4632 5138 4684
rect 5813 4675 5871 4681
rect 5813 4641 5825 4675
rect 5859 4641 5871 4675
rect 5813 4635 5871 4641
rect 4801 4607 4859 4613
rect 4801 4604 4813 4607
rect 4632 4576 4813 4604
rect 4801 4573 4813 4576
rect 4847 4573 4859 4607
rect 4801 4567 4859 4573
rect 5626 4564 5632 4616
rect 5684 4564 5690 4616
rect 4433 4539 4491 4545
rect 4433 4505 4445 4539
rect 4479 4536 4491 4539
rect 4890 4536 4896 4548
rect 4479 4508 4896 4536
rect 4479 4505 4491 4508
rect 4433 4499 4491 4505
rect 4890 4496 4896 4508
rect 4948 4496 4954 4548
rect 5442 4536 5448 4548
rect 5000 4508 5448 4536
rect 4522 4468 4528 4480
rect 4356 4440 4528 4468
rect 4522 4428 4528 4440
rect 4580 4468 4586 4480
rect 4706 4468 4712 4480
rect 4580 4440 4712 4468
rect 4580 4428 4586 4440
rect 4706 4428 4712 4440
rect 4764 4428 4770 4480
rect 5000 4477 5028 4508
rect 5442 4496 5448 4508
rect 5500 4536 5506 4548
rect 5500 4508 5663 4536
rect 5500 4496 5506 4508
rect 4985 4471 5043 4477
rect 4985 4437 4997 4471
rect 5031 4437 5043 4471
rect 4985 4431 5043 4437
rect 5169 4471 5227 4477
rect 5169 4437 5181 4471
rect 5215 4468 5227 4471
rect 5534 4468 5540 4480
rect 5215 4440 5540 4468
rect 5215 4437 5227 4440
rect 5169 4431 5227 4437
rect 5534 4428 5540 4440
rect 5592 4428 5598 4480
rect 5635 4468 5663 4508
rect 5828 4468 5856 4635
rect 6104 4613 6132 4712
rect 6178 4632 6184 4684
rect 6236 4632 6242 4684
rect 7484 4672 7512 4768
rect 6380 4644 7512 4672
rect 8220 4672 8248 4768
rect 8220 4644 8708 4672
rect 6089 4607 6147 4613
rect 6089 4573 6101 4607
rect 6135 4573 6147 4607
rect 6196 4604 6224 4632
rect 6273 4607 6331 4613
rect 6273 4604 6285 4607
rect 6196 4576 6285 4604
rect 6089 4567 6147 4573
rect 6273 4573 6285 4576
rect 6319 4573 6331 4607
rect 6273 4567 6331 4573
rect 6380 4536 6408 4644
rect 6454 4564 6460 4616
rect 6512 4564 6518 4616
rect 7006 4564 7012 4616
rect 7064 4564 7070 4616
rect 7190 4564 7196 4616
rect 7248 4564 7254 4616
rect 7469 4607 7527 4613
rect 7469 4573 7481 4607
rect 7515 4604 7527 4607
rect 7653 4607 7711 4613
rect 7653 4604 7665 4607
rect 7515 4576 7665 4604
rect 7515 4573 7527 4576
rect 7469 4567 7527 4573
rect 7653 4573 7665 4576
rect 7699 4573 7711 4607
rect 7653 4567 7711 4573
rect 8294 4564 8300 4616
rect 8352 4564 8358 4616
rect 8680 4613 8708 4644
rect 8665 4607 8723 4613
rect 8665 4573 8677 4607
rect 8711 4573 8723 4607
rect 8665 4567 8723 4573
rect 5920 4508 6408 4536
rect 6472 4508 7052 4536
rect 5920 4480 5948 4508
rect 5635 4440 5856 4468
rect 5902 4428 5908 4480
rect 5960 4428 5966 4480
rect 5994 4428 6000 4480
rect 6052 4428 6058 4480
rect 6178 4428 6184 4480
rect 6236 4468 6242 4480
rect 6472 4468 6500 4508
rect 6236 4440 6500 4468
rect 6236 4428 6242 4440
rect 6822 4428 6828 4480
rect 6880 4428 6886 4480
rect 7024 4468 7052 4508
rect 7098 4496 7104 4548
rect 7156 4496 7162 4548
rect 7311 4539 7369 4545
rect 7311 4505 7323 4539
rect 7357 4505 7369 4539
rect 7311 4499 7369 4505
rect 7326 4468 7354 4499
rect 8570 4496 8576 4548
rect 8628 4496 8634 4548
rect 7024 4440 7354 4468
rect 1104 4378 9016 4400
rect 1104 4326 2599 4378
rect 2651 4326 2663 4378
rect 2715 4326 2727 4378
rect 2779 4326 2791 4378
rect 2843 4326 2855 4378
rect 2907 4326 4577 4378
rect 4629 4326 4641 4378
rect 4693 4326 4705 4378
rect 4757 4326 4769 4378
rect 4821 4326 4833 4378
rect 4885 4326 6555 4378
rect 6607 4326 6619 4378
rect 6671 4326 6683 4378
rect 6735 4326 6747 4378
rect 6799 4326 6811 4378
rect 6863 4326 8533 4378
rect 8585 4326 8597 4378
rect 8649 4326 8661 4378
rect 8713 4326 8725 4378
rect 8777 4326 8789 4378
rect 8841 4326 9016 4378
rect 1104 4304 9016 4326
rect 1946 4224 1952 4276
rect 2004 4224 2010 4276
rect 3329 4267 3387 4273
rect 3329 4233 3341 4267
rect 3375 4264 3387 4267
rect 3375 4236 4108 4264
rect 3375 4233 3387 4236
rect 3329 4227 3387 4233
rect 1964 4196 1992 4224
rect 2317 4199 2375 4205
rect 2317 4196 2329 4199
rect 1964 4168 2329 4196
rect 2317 4165 2329 4168
rect 2363 4165 2375 4199
rect 3970 4196 3976 4208
rect 2317 4159 2375 4165
rect 2884 4168 3976 4196
rect 1486 4088 1492 4140
rect 1544 4088 1550 4140
rect 1670 4088 1676 4140
rect 1728 4088 1734 4140
rect 1949 4131 2007 4137
rect 1949 4097 1961 4131
rect 1995 4097 2007 4131
rect 1949 4091 2007 4097
rect 2128 4121 2186 4127
rect 1673 3995 1731 4001
rect 1673 3961 1685 3995
rect 1719 3992 1731 3995
rect 1762 3992 1768 4004
rect 1719 3964 1768 3992
rect 1719 3961 1731 3964
rect 1673 3955 1731 3961
rect 1762 3952 1768 3964
rect 1820 3952 1826 4004
rect 1854 3884 1860 3936
rect 1912 3884 1918 3936
rect 1964 3924 1992 4091
rect 2128 4087 2140 4121
rect 2174 4087 2186 4121
rect 2222 4088 2228 4140
rect 2280 4088 2286 4140
rect 2501 4131 2559 4137
rect 2501 4097 2513 4131
rect 2547 4128 2559 4131
rect 2593 4131 2651 4137
rect 2593 4128 2605 4131
rect 2547 4100 2605 4128
rect 2547 4097 2559 4100
rect 2501 4091 2559 4097
rect 2593 4097 2605 4100
rect 2639 4097 2651 4131
rect 2593 4091 2651 4097
rect 2128 4081 2186 4087
rect 2148 3992 2176 4081
rect 2314 4020 2320 4072
rect 2372 4060 2378 4072
rect 2884 4060 2912 4168
rect 3970 4156 3976 4168
rect 4028 4156 4034 4208
rect 2958 4088 2964 4140
rect 3016 4128 3022 4140
rect 3237 4131 3295 4137
rect 3237 4128 3249 4131
rect 3016 4100 3249 4128
rect 3016 4088 3022 4100
rect 3237 4097 3249 4100
rect 3283 4128 3295 4131
rect 3786 4128 3792 4140
rect 3283 4100 3792 4128
rect 3283 4097 3295 4100
rect 3237 4091 3295 4097
rect 3786 4088 3792 4100
rect 3844 4088 3850 4140
rect 2372 4032 2912 4060
rect 3973 4063 4031 4069
rect 2372 4020 2378 4032
rect 3973 4029 3985 4063
rect 4019 4029 4031 4063
rect 4080 4060 4108 4236
rect 4154 4224 4160 4276
rect 4212 4264 4218 4276
rect 5902 4264 5908 4276
rect 4212 4236 5908 4264
rect 4212 4224 4218 4236
rect 5902 4224 5908 4236
rect 5960 4224 5966 4276
rect 6181 4267 6239 4273
rect 6181 4233 6193 4267
rect 6227 4264 6239 4267
rect 7098 4264 7104 4276
rect 6227 4236 7104 4264
rect 6227 4233 6239 4236
rect 6181 4227 6239 4233
rect 7098 4224 7104 4236
rect 7156 4224 7162 4276
rect 8386 4224 8392 4276
rect 8444 4264 8450 4276
rect 8573 4267 8631 4273
rect 8573 4264 8585 4267
rect 8444 4236 8585 4264
rect 8444 4224 8450 4236
rect 8573 4233 8585 4236
rect 8619 4233 8631 4267
rect 8573 4227 8631 4233
rect 4172 4137 4200 4224
rect 5534 4196 5540 4208
rect 5368 4168 5540 4196
rect 4157 4131 4215 4137
rect 4157 4097 4169 4131
rect 4203 4097 4215 4131
rect 4157 4091 4215 4097
rect 4982 4088 4988 4140
rect 5040 4088 5046 4140
rect 5077 4131 5135 4137
rect 5077 4097 5089 4131
rect 5123 4097 5135 4131
rect 5077 4091 5135 4097
rect 4522 4060 4528 4072
rect 4080 4032 4528 4060
rect 3973 4023 4031 4029
rect 2866 3992 2872 4004
rect 2148 3964 2872 3992
rect 2866 3952 2872 3964
rect 2924 3952 2930 4004
rect 3234 3952 3240 4004
rect 3292 3992 3298 4004
rect 3988 3992 4016 4023
rect 4522 4020 4528 4032
rect 4580 4060 4586 4072
rect 5092 4060 5120 4091
rect 4580 4032 5120 4060
rect 4580 4020 4586 4032
rect 4062 3992 4068 4004
rect 3292 3964 4068 3992
rect 3292 3952 3298 3964
rect 4062 3952 4068 3964
rect 4120 3992 4126 4004
rect 5368 3992 5396 4168
rect 5534 4156 5540 4168
rect 5592 4196 5598 4208
rect 5813 4199 5871 4205
rect 5813 4196 5825 4199
rect 5592 4168 5825 4196
rect 5592 4156 5598 4168
rect 5813 4165 5825 4168
rect 5859 4165 5871 4199
rect 5813 4159 5871 4165
rect 6043 4165 6101 4171
rect 5445 4131 5503 4137
rect 5445 4097 5457 4131
rect 5491 4128 5503 4131
rect 5491 4100 5580 4128
rect 5491 4097 5503 4100
rect 5445 4091 5503 4097
rect 4120 3964 5396 3992
rect 4120 3952 4126 3964
rect 5552 3936 5580 4100
rect 5626 4088 5632 4140
rect 5684 4128 5690 4140
rect 6043 4131 6055 4165
rect 6089 4131 6101 4165
rect 6472 4168 7604 4196
rect 6043 4128 6101 4131
rect 6270 4128 6276 4140
rect 5684 4100 6276 4128
rect 5684 4088 5690 4100
rect 6270 4088 6276 4100
rect 6328 4088 6334 4140
rect 6365 4131 6423 4137
rect 6365 4097 6377 4131
rect 6411 4128 6423 4131
rect 6472 4128 6500 4168
rect 7576 4140 7604 4168
rect 6411 4100 6500 4128
rect 6549 4131 6607 4137
rect 6411 4097 6423 4100
rect 6365 4091 6423 4097
rect 6549 4097 6561 4131
rect 6595 4097 6607 4131
rect 6549 4091 6607 4097
rect 6641 4131 6699 4137
rect 6641 4097 6653 4131
rect 6687 4128 6699 4131
rect 6733 4131 6791 4137
rect 6687 4097 6700 4128
rect 6641 4091 6700 4097
rect 6733 4097 6745 4131
rect 6779 4128 6791 4131
rect 6822 4128 6828 4140
rect 6779 4100 6828 4128
rect 6779 4097 6791 4100
rect 6733 4091 6791 4097
rect 6178 4060 6184 4072
rect 5644 4032 6184 4060
rect 5644 3936 5672 4032
rect 6178 4020 6184 4032
rect 6236 4060 6242 4072
rect 6564 4060 6592 4091
rect 6236 4032 6592 4060
rect 6236 4020 6242 4032
rect 2406 3924 2412 3936
rect 1964 3896 2412 3924
rect 2406 3884 2412 3896
rect 2464 3884 2470 3936
rect 2498 3884 2504 3936
rect 2556 3884 2562 3936
rect 5534 3884 5540 3936
rect 5592 3884 5598 3936
rect 5626 3884 5632 3936
rect 5684 3884 5690 3936
rect 5997 3927 6055 3933
rect 5997 3893 6009 3927
rect 6043 3924 6055 3927
rect 6362 3924 6368 3936
rect 6043 3896 6368 3924
rect 6043 3893 6055 3896
rect 5997 3887 6055 3893
rect 6362 3884 6368 3896
rect 6420 3884 6426 3936
rect 6672 3924 6700 4091
rect 6822 4088 6828 4100
rect 6880 4088 6886 4140
rect 7009 4131 7067 4137
rect 7009 4097 7021 4131
rect 7055 4097 7067 4131
rect 7009 4091 7067 4097
rect 7024 4060 7052 4091
rect 7098 4088 7104 4140
rect 7156 4128 7162 4140
rect 7265 4131 7323 4137
rect 7265 4128 7277 4131
rect 7156 4100 7277 4128
rect 7156 4088 7162 4100
rect 7265 4097 7277 4100
rect 7311 4097 7323 4131
rect 7265 4091 7323 4097
rect 7558 4088 7564 4140
rect 7616 4088 7622 4140
rect 8665 4131 8723 4137
rect 8665 4097 8677 4131
rect 8711 4128 8723 4131
rect 8938 4128 8944 4140
rect 8711 4100 8944 4128
rect 8711 4097 8723 4100
rect 8665 4091 8723 4097
rect 8938 4088 8944 4100
rect 8996 4088 9002 4140
rect 6748 4032 7052 4060
rect 6748 4004 6776 4032
rect 8294 4020 8300 4072
rect 8352 4020 8358 4072
rect 6730 3952 6736 4004
rect 6788 3952 6794 4004
rect 6917 3995 6975 4001
rect 6917 3961 6929 3995
rect 6963 3992 6975 3995
rect 7006 3992 7012 4004
rect 6963 3964 7012 3992
rect 6963 3961 6975 3964
rect 6917 3955 6975 3961
rect 7006 3952 7012 3964
rect 7064 3952 7070 4004
rect 8312 3992 8340 4020
rect 8389 3995 8447 4001
rect 8389 3992 8401 3995
rect 8312 3964 8401 3992
rect 8389 3961 8401 3964
rect 8435 3961 8447 3995
rect 8389 3955 8447 3961
rect 7190 3924 7196 3936
rect 6672 3896 7196 3924
rect 7190 3884 7196 3896
rect 7248 3884 7254 3936
rect 1104 3834 9016 3856
rect 1104 3782 1939 3834
rect 1991 3782 2003 3834
rect 2055 3782 2067 3834
rect 2119 3782 2131 3834
rect 2183 3782 2195 3834
rect 2247 3782 3917 3834
rect 3969 3782 3981 3834
rect 4033 3782 4045 3834
rect 4097 3782 4109 3834
rect 4161 3782 4173 3834
rect 4225 3782 5895 3834
rect 5947 3782 5959 3834
rect 6011 3782 6023 3834
rect 6075 3782 6087 3834
rect 6139 3782 6151 3834
rect 6203 3782 7873 3834
rect 7925 3782 7937 3834
rect 7989 3782 8001 3834
rect 8053 3782 8065 3834
rect 8117 3782 8129 3834
rect 8181 3782 9016 3834
rect 1104 3760 9016 3782
rect 2498 3680 2504 3732
rect 2556 3680 2562 3732
rect 2866 3680 2872 3732
rect 2924 3680 2930 3732
rect 3418 3720 3424 3732
rect 3252 3692 3424 3720
rect 1394 3544 1400 3596
rect 1452 3544 1458 3596
rect 1664 3519 1722 3525
rect 1664 3485 1676 3519
rect 1710 3516 1722 3519
rect 2516 3516 2544 3680
rect 2777 3655 2835 3661
rect 2777 3621 2789 3655
rect 2823 3652 2835 3655
rect 3252 3652 3280 3692
rect 3418 3680 3424 3692
rect 3476 3680 3482 3732
rect 3602 3720 3608 3732
rect 3600 3680 3608 3720
rect 3660 3680 3666 3732
rect 3694 3680 3700 3732
rect 3752 3720 3758 3732
rect 4341 3723 4399 3729
rect 4341 3720 4353 3723
rect 3752 3692 4353 3720
rect 3752 3680 3758 3692
rect 4341 3689 4353 3692
rect 4387 3689 4399 3723
rect 4341 3683 4399 3689
rect 4614 3680 4620 3732
rect 4672 3720 4678 3732
rect 5534 3720 5540 3732
rect 4672 3692 5540 3720
rect 4672 3680 4678 3692
rect 5534 3680 5540 3692
rect 5592 3720 5598 3732
rect 6825 3723 6883 3729
rect 6825 3720 6837 3723
rect 5592 3692 6837 3720
rect 5592 3680 5598 3692
rect 6825 3689 6837 3692
rect 6871 3689 6883 3723
rect 6825 3683 6883 3689
rect 7193 3723 7251 3729
rect 7193 3689 7205 3723
rect 7239 3720 7251 3723
rect 7466 3720 7472 3732
rect 7239 3692 7472 3720
rect 7239 3689 7251 3692
rect 7193 3683 7251 3689
rect 7466 3680 7472 3692
rect 7524 3680 7530 3732
rect 2823 3624 3280 3652
rect 2823 3621 2835 3624
rect 2777 3615 2835 3621
rect 3326 3612 3332 3664
rect 3384 3612 3390 3664
rect 2958 3584 2964 3596
rect 2884 3556 2964 3584
rect 2884 3525 2912 3556
rect 2958 3544 2964 3556
rect 3016 3544 3022 3596
rect 3050 3544 3056 3596
rect 3108 3544 3114 3596
rect 3600 3584 3628 3680
rect 5166 3612 5172 3664
rect 5224 3612 5230 3664
rect 6730 3584 6736 3596
rect 3160 3556 3628 3584
rect 3160 3525 3188 3556
rect 1710 3488 2544 3516
rect 2869 3519 2927 3525
rect 1710 3485 1722 3488
rect 1664 3479 1722 3485
rect 2869 3485 2881 3519
rect 2915 3485 2927 3519
rect 2869 3479 2927 3485
rect 3145 3519 3203 3525
rect 3145 3485 3157 3519
rect 3191 3485 3203 3519
rect 3145 3479 3203 3485
rect 3234 3476 3240 3528
rect 3292 3476 3298 3528
rect 3600 3525 3628 3556
rect 3804 3556 4568 3584
rect 3804 3525 3832 3556
rect 4540 3528 4568 3556
rect 6472 3556 6736 3584
rect 3600 3519 3663 3525
rect 3600 3488 3617 3519
rect 3605 3485 3617 3488
rect 3651 3485 3663 3519
rect 3605 3479 3663 3485
rect 3789 3519 3847 3525
rect 3789 3485 3801 3519
rect 3835 3485 3847 3519
rect 3789 3479 3847 3485
rect 3878 3476 3884 3528
rect 3936 3476 3942 3528
rect 4157 3519 4215 3525
rect 4157 3485 4169 3519
rect 4203 3485 4215 3519
rect 4157 3479 4215 3485
rect 4249 3519 4307 3525
rect 4249 3485 4261 3519
rect 4295 3516 4307 3519
rect 4430 3516 4436 3528
rect 4295 3488 4436 3516
rect 4295 3485 4307 3488
rect 4249 3479 4307 3485
rect 3329 3451 3387 3457
rect 3329 3417 3341 3451
rect 3375 3448 3387 3451
rect 3418 3448 3424 3460
rect 3375 3420 3424 3448
rect 3375 3417 3387 3420
rect 3329 3411 3387 3417
rect 3418 3408 3424 3420
rect 3476 3448 3482 3460
rect 3896 3448 3924 3476
rect 3476 3420 3924 3448
rect 3476 3408 3482 3420
rect 3050 3340 3056 3392
rect 3108 3380 3114 3392
rect 3513 3383 3571 3389
rect 3513 3380 3525 3383
rect 3108 3352 3525 3380
rect 3108 3340 3114 3352
rect 3513 3349 3525 3352
rect 3559 3380 3571 3383
rect 3786 3380 3792 3392
rect 3559 3352 3792 3380
rect 3559 3349 3571 3352
rect 3513 3343 3571 3349
rect 3786 3340 3792 3352
rect 3844 3340 3850 3392
rect 3878 3340 3884 3392
rect 3936 3340 3942 3392
rect 3970 3340 3976 3392
rect 4028 3340 4034 3392
rect 4062 3340 4068 3392
rect 4120 3340 4126 3392
rect 4172 3380 4200 3479
rect 4430 3476 4436 3488
rect 4488 3476 4494 3528
rect 4522 3476 4528 3528
rect 4580 3476 4586 3528
rect 4614 3476 4620 3528
rect 4672 3476 4678 3528
rect 4709 3519 4767 3525
rect 4709 3485 4721 3519
rect 4755 3516 4767 3519
rect 4982 3516 4988 3528
rect 4755 3488 4988 3516
rect 4755 3485 4767 3488
rect 4709 3479 4767 3485
rect 4982 3476 4988 3488
rect 5040 3476 5046 3528
rect 5077 3519 5135 3525
rect 5077 3485 5089 3519
rect 5123 3516 5135 3519
rect 5166 3516 5172 3528
rect 5123 3488 5172 3516
rect 5123 3485 5135 3488
rect 5077 3479 5135 3485
rect 5166 3476 5172 3488
rect 5224 3476 5230 3528
rect 5258 3476 5264 3528
rect 5316 3516 5322 3528
rect 5353 3519 5411 3525
rect 5353 3516 5365 3519
rect 5316 3488 5365 3516
rect 5316 3476 5322 3488
rect 5353 3485 5365 3488
rect 5399 3516 5411 3519
rect 6472 3516 6500 3556
rect 6730 3544 6736 3556
rect 6788 3584 6794 3596
rect 7285 3587 7343 3593
rect 7285 3584 7297 3587
rect 6788 3556 7297 3584
rect 6788 3544 6794 3556
rect 7285 3553 7297 3556
rect 7331 3553 7343 3587
rect 7285 3547 7343 3553
rect 7009 3519 7067 3525
rect 7009 3516 7021 3519
rect 5399 3488 6500 3516
rect 6564 3488 7021 3516
rect 5399 3485 5411 3488
rect 5353 3479 5411 3485
rect 4448 3448 4476 3476
rect 5620 3451 5678 3457
rect 4448 3420 5580 3448
rect 4614 3380 4620 3392
rect 4172 3352 4620 3380
rect 4614 3340 4620 3352
rect 4672 3340 4678 3392
rect 4982 3340 4988 3392
rect 5040 3340 5046 3392
rect 5552 3380 5580 3420
rect 5620 3417 5632 3451
rect 5666 3448 5678 3451
rect 6270 3448 6276 3460
rect 5666 3420 6276 3448
rect 5666 3417 5678 3420
rect 5620 3411 5678 3417
rect 6270 3408 6276 3420
rect 6328 3408 6334 3460
rect 6564 3380 6592 3488
rect 7009 3485 7021 3488
rect 7055 3485 7067 3519
rect 7009 3479 7067 3485
rect 7098 3476 7104 3528
rect 7156 3476 7162 3528
rect 7193 3519 7251 3525
rect 7193 3485 7205 3519
rect 7239 3516 7251 3519
rect 7541 3519 7599 3525
rect 7541 3516 7553 3519
rect 7239 3488 7328 3516
rect 7239 3485 7251 3488
rect 7193 3479 7251 3485
rect 5552 3352 6592 3380
rect 6733 3383 6791 3389
rect 6733 3349 6745 3383
rect 6779 3380 6791 3383
rect 7006 3380 7012 3392
rect 6779 3352 7012 3380
rect 6779 3349 6791 3352
rect 6733 3343 6791 3349
rect 7006 3340 7012 3352
rect 7064 3340 7070 3392
rect 7116 3380 7144 3476
rect 7300 3460 7328 3488
rect 7392 3488 7553 3516
rect 7282 3408 7288 3460
rect 7340 3408 7346 3460
rect 7392 3380 7420 3488
rect 7541 3485 7553 3488
rect 7587 3485 7599 3519
rect 7541 3479 7599 3485
rect 7116 3352 7420 3380
rect 8665 3383 8723 3389
rect 8665 3349 8677 3383
rect 8711 3380 8723 3383
rect 8711 3352 9076 3380
rect 8711 3349 8723 3352
rect 8665 3343 8723 3349
rect 1104 3290 9016 3312
rect 1104 3238 2599 3290
rect 2651 3238 2663 3290
rect 2715 3238 2727 3290
rect 2779 3238 2791 3290
rect 2843 3238 2855 3290
rect 2907 3238 4577 3290
rect 4629 3238 4641 3290
rect 4693 3238 4705 3290
rect 4757 3238 4769 3290
rect 4821 3238 4833 3290
rect 4885 3238 6555 3290
rect 6607 3238 6619 3290
rect 6671 3238 6683 3290
rect 6735 3238 6747 3290
rect 6799 3238 6811 3290
rect 6863 3238 8533 3290
rect 8585 3238 8597 3290
rect 8649 3238 8661 3290
rect 8713 3238 8725 3290
rect 8777 3238 8789 3290
rect 8841 3238 9016 3290
rect 1104 3216 9016 3238
rect 1394 3136 1400 3188
rect 1452 3136 1458 3188
rect 1854 3136 1860 3188
rect 1912 3176 1918 3188
rect 1912 3148 4108 3176
rect 1912 3136 1918 3148
rect 1412 3108 1440 3136
rect 2593 3111 2651 3117
rect 2593 3108 2605 3111
rect 1412 3080 2605 3108
rect 2593 3077 2605 3080
rect 2639 3108 2651 3111
rect 2774 3108 2780 3120
rect 2639 3080 2780 3108
rect 2639 3077 2651 3080
rect 2593 3071 2651 3077
rect 2774 3068 2780 3080
rect 2832 3068 2838 3120
rect 1762 3000 1768 3052
rect 1820 3049 1826 3052
rect 1820 3043 1841 3049
rect 1829 3009 1841 3043
rect 1820 3003 1841 3009
rect 1820 3000 1826 3003
rect 2038 3000 2044 3052
rect 2096 3000 2102 3052
rect 2317 3043 2375 3049
rect 2317 3009 2329 3043
rect 2363 3009 2375 3043
rect 2317 3003 2375 3009
rect 2501 3043 2559 3049
rect 2501 3009 2513 3043
rect 2547 3040 2559 3043
rect 3602 3040 3608 3052
rect 2547 3012 3608 3040
rect 2547 3009 2559 3012
rect 2501 3003 2559 3009
rect 2332 2904 2360 3003
rect 3602 3000 3608 3012
rect 3660 3000 3666 3052
rect 4080 3040 4108 3148
rect 4154 3136 4160 3188
rect 4212 3176 4218 3188
rect 4890 3176 4896 3188
rect 4212 3148 4896 3176
rect 4212 3136 4218 3148
rect 4890 3136 4896 3148
rect 4948 3136 4954 3188
rect 4982 3136 4988 3188
rect 5040 3136 5046 3188
rect 5626 3176 5632 3188
rect 5460 3148 5632 3176
rect 4338 3068 4344 3120
rect 4396 3068 4402 3120
rect 5000 3108 5028 3136
rect 5169 3111 5227 3117
rect 5169 3108 5181 3111
rect 5000 3080 5181 3108
rect 5169 3077 5181 3080
rect 5215 3077 5227 3111
rect 5169 3071 5227 3077
rect 5460 3049 5488 3148
rect 5626 3136 5632 3148
rect 5684 3176 5690 3188
rect 6730 3176 6736 3188
rect 5684 3148 6736 3176
rect 5684 3136 5690 3148
rect 6730 3136 6736 3148
rect 6788 3136 6794 3188
rect 6825 3179 6883 3185
rect 6825 3145 6837 3179
rect 6871 3176 6883 3179
rect 6914 3176 6920 3188
rect 6871 3148 6920 3176
rect 6871 3145 6883 3148
rect 6825 3139 6883 3145
rect 6914 3136 6920 3148
rect 6972 3136 6978 3188
rect 7006 3136 7012 3188
rect 7064 3176 7070 3188
rect 7064 3148 7512 3176
rect 7064 3136 7070 3148
rect 5534 3068 5540 3120
rect 5592 3108 5598 3120
rect 6457 3111 6515 3117
rect 6457 3108 6469 3111
rect 5592 3080 6469 3108
rect 5592 3068 5598 3080
rect 6457 3077 6469 3080
rect 6503 3077 6515 3111
rect 7374 3108 7380 3120
rect 6457 3071 6515 3077
rect 6687 3077 6745 3083
rect 5353 3043 5411 3049
rect 5353 3040 5365 3043
rect 4080 3012 5365 3040
rect 5353 3009 5365 3012
rect 5399 3009 5411 3043
rect 5353 3003 5411 3009
rect 5445 3043 5503 3049
rect 5445 3009 5457 3043
rect 5491 3009 5503 3043
rect 5445 3003 5503 3009
rect 5552 3012 5856 3040
rect 2409 2975 2467 2981
rect 2409 2941 2421 2975
rect 2455 2972 2467 2975
rect 2455 2944 4476 2972
rect 2455 2941 2467 2944
rect 2409 2935 2467 2941
rect 3234 2904 3240 2916
rect 2332 2876 3240 2904
rect 3234 2864 3240 2876
rect 3292 2864 3298 2916
rect 4448 2904 4476 2944
rect 4982 2932 4988 2984
rect 5040 2972 5046 2984
rect 5552 2972 5580 3012
rect 5040 2944 5580 2972
rect 5040 2932 5046 2944
rect 5626 2932 5632 2984
rect 5684 2932 5690 2984
rect 5828 2972 5856 3012
rect 5902 3000 5908 3052
rect 5960 3040 5966 3052
rect 6687 3043 6699 3077
rect 6733 3043 6745 3077
rect 6932 3080 7380 3108
rect 6932 3052 6960 3080
rect 7374 3068 7380 3080
rect 7432 3068 7438 3120
rect 6687 3040 6745 3043
rect 5960 3037 6745 3040
rect 5960 3012 6730 3037
rect 5960 3000 5966 3012
rect 6914 3000 6920 3052
rect 6972 3000 6978 3052
rect 7190 3040 7196 3052
rect 7024 3012 7196 3040
rect 7024 2972 7052 3012
rect 7190 3000 7196 3012
rect 7248 3000 7254 3052
rect 7484 2972 7512 3148
rect 8018 3136 8024 3188
rect 8076 3136 8082 3188
rect 8205 3179 8263 3185
rect 8205 3145 8217 3179
rect 8251 3176 8263 3179
rect 8294 3176 8300 3188
rect 8251 3148 8300 3176
rect 8251 3145 8263 3148
rect 8205 3139 8263 3145
rect 7561 3043 7619 3049
rect 7561 3009 7573 3043
rect 7607 3040 7619 3043
rect 7742 3040 7748 3052
rect 7607 3012 7748 3040
rect 7607 3009 7619 3012
rect 7561 3003 7619 3009
rect 7742 3000 7748 3012
rect 7800 3040 7806 3052
rect 8220 3040 8248 3139
rect 8294 3136 8300 3148
rect 8352 3136 8358 3188
rect 9048 3176 9076 3352
rect 8680 3148 9076 3176
rect 7800 3012 8248 3040
rect 8297 3043 8355 3049
rect 7800 3000 7806 3012
rect 8297 3009 8309 3043
rect 8343 3009 8355 3043
rect 8297 3003 8355 3009
rect 8389 3043 8447 3049
rect 8389 3009 8401 3043
rect 8435 3040 8447 3043
rect 8680 3040 8708 3148
rect 8435 3012 8708 3040
rect 8435 3009 8447 3012
rect 8389 3003 8447 3009
rect 7929 2975 7987 2981
rect 7929 2972 7941 2975
rect 5828 2944 7144 2972
rect 7484 2944 7941 2972
rect 5810 2904 5816 2916
rect 4448 2876 5816 2904
rect 5810 2864 5816 2876
rect 5868 2864 5874 2916
rect 7006 2904 7012 2916
rect 6656 2876 7012 2904
rect 14 2796 20 2848
rect 72 2836 78 2848
rect 1489 2839 1547 2845
rect 1489 2836 1501 2839
rect 72 2808 1501 2836
rect 72 2796 78 2808
rect 1489 2805 1501 2808
rect 1535 2805 1547 2839
rect 1489 2799 1547 2805
rect 2225 2839 2283 2845
rect 2225 2805 2237 2839
rect 2271 2836 2283 2839
rect 2314 2836 2320 2848
rect 2271 2808 2320 2836
rect 2271 2805 2283 2808
rect 2225 2799 2283 2805
rect 2314 2796 2320 2808
rect 2372 2796 2378 2848
rect 2590 2796 2596 2848
rect 2648 2836 2654 2848
rect 4433 2839 4491 2845
rect 4433 2836 4445 2839
rect 2648 2808 4445 2836
rect 2648 2796 2654 2808
rect 4433 2805 4445 2808
rect 4479 2805 4491 2839
rect 4433 2799 4491 2805
rect 5166 2796 5172 2848
rect 5224 2796 5230 2848
rect 6181 2839 6239 2845
rect 6181 2805 6193 2839
rect 6227 2836 6239 2839
rect 6362 2836 6368 2848
rect 6227 2808 6368 2836
rect 6227 2805 6239 2808
rect 6181 2799 6239 2805
rect 6362 2796 6368 2808
rect 6420 2796 6426 2848
rect 6656 2845 6684 2876
rect 7006 2864 7012 2876
rect 7064 2864 7070 2916
rect 7116 2904 7144 2944
rect 7929 2941 7941 2944
rect 7975 2972 7987 2975
rect 8312 2972 8340 3003
rect 8478 2972 8484 2984
rect 7975 2944 8484 2972
rect 7975 2941 7987 2944
rect 7929 2935 7987 2941
rect 8478 2932 8484 2944
rect 8536 2932 8542 2984
rect 8573 2907 8631 2913
rect 8573 2904 8585 2907
rect 7116 2876 8585 2904
rect 8573 2873 8585 2876
rect 8619 2873 8631 2907
rect 8573 2867 8631 2873
rect 6641 2839 6699 2845
rect 6641 2805 6653 2839
rect 6687 2805 6699 2839
rect 6641 2799 6699 2805
rect 6822 2796 6828 2848
rect 6880 2836 6886 2848
rect 7469 2839 7527 2845
rect 7469 2836 7481 2839
rect 6880 2808 7481 2836
rect 6880 2796 6886 2808
rect 7469 2805 7481 2808
rect 7515 2805 7527 2839
rect 7469 2799 7527 2805
rect 7650 2796 7656 2848
rect 7708 2836 7714 2848
rect 8294 2836 8300 2848
rect 7708 2808 8300 2836
rect 7708 2796 7714 2808
rect 8294 2796 8300 2808
rect 8352 2836 8358 2848
rect 8680 2836 8708 3012
rect 8352 2808 8708 2836
rect 8352 2796 8358 2808
rect 1104 2746 9016 2768
rect 1104 2694 1939 2746
rect 1991 2694 2003 2746
rect 2055 2694 2067 2746
rect 2119 2694 2131 2746
rect 2183 2694 2195 2746
rect 2247 2694 3917 2746
rect 3969 2694 3981 2746
rect 4033 2694 4045 2746
rect 4097 2694 4109 2746
rect 4161 2694 4173 2746
rect 4225 2694 5895 2746
rect 5947 2694 5959 2746
rect 6011 2694 6023 2746
rect 6075 2694 6087 2746
rect 6139 2694 6151 2746
rect 6203 2694 7873 2746
rect 7925 2694 7937 2746
rect 7989 2694 8001 2746
rect 8053 2694 8065 2746
rect 8117 2694 8129 2746
rect 8181 2694 9016 2746
rect 1104 2672 9016 2694
rect 1397 2635 1455 2641
rect 1397 2601 1409 2635
rect 1443 2632 1455 2635
rect 1762 2632 1768 2644
rect 1443 2604 1768 2632
rect 1443 2601 1455 2604
rect 1397 2595 1455 2601
rect 1762 2592 1768 2604
rect 1820 2632 1826 2644
rect 2498 2632 2504 2644
rect 1820 2604 2504 2632
rect 1820 2592 1826 2604
rect 2498 2592 2504 2604
rect 2556 2592 2562 2644
rect 2774 2592 2780 2644
rect 2832 2592 2838 2644
rect 3602 2592 3608 2644
rect 3660 2632 3666 2644
rect 3881 2635 3939 2641
rect 3881 2632 3893 2635
rect 3660 2604 3893 2632
rect 3660 2592 3666 2604
rect 3881 2601 3893 2604
rect 3927 2632 3939 2635
rect 4982 2632 4988 2644
rect 3927 2604 4988 2632
rect 3927 2601 3939 2604
rect 3881 2595 3939 2601
rect 4982 2592 4988 2604
rect 5040 2592 5046 2644
rect 5626 2592 5632 2644
rect 5684 2632 5690 2644
rect 5902 2632 5908 2644
rect 5684 2604 5908 2632
rect 5684 2592 5690 2604
rect 5902 2592 5908 2604
rect 5960 2592 5966 2644
rect 6270 2592 6276 2644
rect 6328 2632 6334 2644
rect 6641 2635 6699 2641
rect 6641 2632 6653 2635
rect 6328 2604 6653 2632
rect 6328 2592 6334 2604
rect 6641 2601 6653 2604
rect 6687 2601 6699 2635
rect 6641 2595 6699 2601
rect 7006 2592 7012 2644
rect 7064 2592 7070 2644
rect 7116 2604 8616 2632
rect 2792 2564 2820 2592
rect 6454 2564 6460 2576
rect 2792 2536 4200 2564
rect 2792 2505 2820 2536
rect 2777 2499 2835 2505
rect 2777 2465 2789 2499
rect 2823 2465 2835 2499
rect 3053 2499 3111 2505
rect 3053 2496 3065 2499
rect 2777 2459 2835 2465
rect 2884 2468 3065 2496
rect 2521 2431 2579 2437
rect 2521 2397 2533 2431
rect 2567 2428 2579 2431
rect 2884 2428 2912 2468
rect 3053 2465 3065 2468
rect 3099 2465 3111 2499
rect 3053 2459 3111 2465
rect 3234 2456 3240 2508
rect 3292 2456 3298 2508
rect 3528 2468 3740 2496
rect 2567 2400 2912 2428
rect 2956 2431 3014 2437
rect 2567 2397 2579 2400
rect 2521 2391 2579 2397
rect 2956 2397 2968 2431
rect 3002 2428 3014 2431
rect 3252 2428 3280 2456
rect 3002 2400 3280 2428
rect 3002 2397 3014 2400
rect 2956 2391 3014 2397
rect 3326 2388 3332 2440
rect 3384 2388 3390 2440
rect 3418 2388 3424 2440
rect 3476 2388 3482 2440
rect 3050 2320 3056 2372
rect 3108 2320 3114 2372
rect 3145 2363 3203 2369
rect 3145 2329 3157 2363
rect 3191 2360 3203 2363
rect 3528 2360 3556 2468
rect 3605 2431 3663 2437
rect 3605 2397 3617 2431
rect 3651 2397 3663 2431
rect 3605 2391 3663 2397
rect 3191 2332 3556 2360
rect 3191 2329 3203 2332
rect 3145 2323 3203 2329
rect 3510 2252 3516 2304
rect 3568 2252 3574 2304
rect 3620 2292 3648 2391
rect 3712 2360 3740 2468
rect 4172 2428 4200 2536
rect 5736 2536 6460 2564
rect 5258 2428 5264 2440
rect 4172 2400 5264 2428
rect 5258 2388 5264 2400
rect 5316 2388 5322 2440
rect 5534 2388 5540 2440
rect 5592 2388 5598 2440
rect 5626 2388 5632 2440
rect 5684 2428 5690 2440
rect 5736 2437 5764 2536
rect 6454 2524 6460 2536
rect 6512 2564 6518 2576
rect 6822 2564 6828 2576
rect 6512 2536 6828 2564
rect 6512 2524 6518 2536
rect 6822 2524 6828 2536
rect 6880 2524 6886 2576
rect 6362 2456 6368 2508
rect 6420 2456 6426 2508
rect 7116 2496 7144 2604
rect 7650 2524 7656 2576
rect 7708 2524 7714 2576
rect 8294 2564 8300 2576
rect 8220 2536 8300 2564
rect 6672 2468 7144 2496
rect 5721 2431 5779 2437
rect 5721 2428 5733 2431
rect 5684 2400 5733 2428
rect 5684 2388 5690 2400
rect 5721 2397 5733 2400
rect 5767 2397 5779 2431
rect 5721 2391 5779 2397
rect 5810 2388 5816 2440
rect 5868 2388 5874 2440
rect 5902 2388 5908 2440
rect 5960 2428 5966 2440
rect 6672 2428 6700 2468
rect 5960 2400 6700 2428
rect 5960 2388 5966 2400
rect 6730 2388 6736 2440
rect 6788 2388 6794 2440
rect 6917 2431 6975 2437
rect 6917 2397 6929 2431
rect 6963 2397 6975 2431
rect 6917 2391 6975 2397
rect 4246 2360 4252 2372
rect 3712 2332 4252 2360
rect 4246 2320 4252 2332
rect 4304 2320 4310 2372
rect 5016 2363 5074 2369
rect 5016 2329 5028 2363
rect 5062 2360 5074 2363
rect 5166 2360 5172 2372
rect 5062 2332 5172 2360
rect 5062 2329 5074 2332
rect 5016 2323 5074 2329
rect 5166 2320 5172 2332
rect 5224 2320 5230 2372
rect 5552 2292 5580 2388
rect 6181 2363 6239 2369
rect 6181 2329 6193 2363
rect 6227 2360 6239 2363
rect 6932 2360 6960 2391
rect 7190 2388 7196 2440
rect 7248 2388 7254 2440
rect 7668 2437 7696 2524
rect 8113 2499 8171 2505
rect 8113 2496 8125 2499
rect 7760 2468 8125 2496
rect 7760 2437 7788 2468
rect 8113 2465 8125 2468
rect 8159 2465 8171 2499
rect 8113 2459 8171 2465
rect 7377 2431 7435 2437
rect 7377 2397 7389 2431
rect 7423 2428 7435 2431
rect 7653 2431 7711 2437
rect 7653 2428 7665 2431
rect 7423 2400 7665 2428
rect 7423 2397 7435 2400
rect 7377 2391 7435 2397
rect 7653 2397 7665 2400
rect 7699 2397 7711 2431
rect 7653 2391 7711 2397
rect 7745 2431 7803 2437
rect 7745 2397 7757 2431
rect 7791 2397 7803 2431
rect 7745 2391 7803 2397
rect 6227 2332 6960 2360
rect 7208 2360 7236 2388
rect 7760 2360 7788 2391
rect 7926 2388 7932 2440
rect 7984 2388 7990 2440
rect 8220 2437 8248 2536
rect 8294 2524 8300 2536
rect 8352 2524 8358 2576
rect 8478 2524 8484 2576
rect 8536 2524 8542 2576
rect 8205 2431 8263 2437
rect 8205 2397 8217 2431
rect 8251 2397 8263 2431
rect 8205 2391 8263 2397
rect 8297 2431 8355 2437
rect 8297 2397 8309 2431
rect 8343 2428 8355 2431
rect 8389 2431 8447 2437
rect 8389 2428 8401 2431
rect 8343 2400 8401 2428
rect 8343 2397 8355 2400
rect 8297 2391 8355 2397
rect 8389 2397 8401 2400
rect 8435 2428 8447 2431
rect 8496 2428 8524 2524
rect 8435 2400 8524 2428
rect 8435 2397 8447 2400
rect 8389 2391 8447 2397
rect 7208 2332 7788 2360
rect 8481 2363 8539 2369
rect 6227 2329 6239 2332
rect 6181 2323 6239 2329
rect 8481 2329 8493 2363
rect 8527 2360 8539 2363
rect 8588 2360 8616 2604
rect 8527 2332 8616 2360
rect 8527 2329 8539 2332
rect 8481 2323 8539 2329
rect 3620 2264 5580 2292
rect 6454 2252 6460 2304
rect 6512 2252 6518 2304
rect 7466 2252 7472 2304
rect 7524 2252 7530 2304
rect 8018 2252 8024 2304
rect 8076 2252 8082 2304
rect 1104 2202 9016 2224
rect 1104 2150 2599 2202
rect 2651 2150 2663 2202
rect 2715 2150 2727 2202
rect 2779 2150 2791 2202
rect 2843 2150 2855 2202
rect 2907 2150 4577 2202
rect 4629 2150 4641 2202
rect 4693 2150 4705 2202
rect 4757 2150 4769 2202
rect 4821 2150 4833 2202
rect 4885 2150 6555 2202
rect 6607 2150 6619 2202
rect 6671 2150 6683 2202
rect 6735 2150 6747 2202
rect 6799 2150 6811 2202
rect 6863 2150 8533 2202
rect 8585 2150 8597 2202
rect 8649 2150 8661 2202
rect 8713 2150 8725 2202
rect 8777 2150 8789 2202
rect 8841 2150 9016 2202
rect 1104 2128 9016 2150
rect 8018 2088 8024 2100
rect 2746 2060 8024 2088
rect 1578 1844 1584 1896
rect 1636 1844 1642 1896
rect 1596 1816 1624 1844
rect 2746 1816 2774 2060
rect 8018 2048 8024 2060
rect 8076 2048 8082 2100
rect 3050 1980 3056 2032
rect 3108 2020 3114 2032
rect 5350 2020 5356 2032
rect 3108 1992 5356 2020
rect 3108 1980 3114 1992
rect 5350 1980 5356 1992
rect 5408 1980 5414 2032
rect 5718 1980 5724 2032
rect 5776 1980 5782 2032
rect 3510 1912 3516 1964
rect 3568 1952 3574 1964
rect 5736 1952 5764 1980
rect 3568 1924 5764 1952
rect 3568 1912 3574 1924
rect 3786 1844 3792 1896
rect 3844 1884 3850 1896
rect 6454 1884 6460 1896
rect 3844 1856 6460 1884
rect 3844 1844 3850 1856
rect 6454 1844 6460 1856
rect 6512 1844 6518 1896
rect 1596 1788 2774 1816
rect 3694 1708 3700 1760
rect 3752 1748 3758 1760
rect 7466 1748 7472 1760
rect 3752 1720 7472 1748
rect 3752 1708 3758 1720
rect 7466 1708 7472 1720
rect 7524 1708 7530 1760
<< via1 >>
rect 2599 9766 2651 9818
rect 2663 9766 2715 9818
rect 2727 9766 2779 9818
rect 2791 9766 2843 9818
rect 2855 9766 2907 9818
rect 4577 9766 4629 9818
rect 4641 9766 4693 9818
rect 4705 9766 4757 9818
rect 4769 9766 4821 9818
rect 4833 9766 4885 9818
rect 6555 9766 6607 9818
rect 6619 9766 6671 9818
rect 6683 9766 6735 9818
rect 6747 9766 6799 9818
rect 6811 9766 6863 9818
rect 8533 9766 8585 9818
rect 8597 9766 8649 9818
rect 8661 9766 8713 9818
rect 8725 9766 8777 9818
rect 8789 9766 8841 9818
rect 2688 9664 2740 9716
rect 2044 9596 2096 9648
rect 1676 9460 1728 9512
rect 1860 9324 1912 9376
rect 2044 9503 2096 9512
rect 2044 9469 2053 9503
rect 2053 9469 2087 9503
rect 2087 9469 2096 9503
rect 2044 9460 2096 9469
rect 2320 9460 2372 9512
rect 2412 9460 2464 9512
rect 3332 9571 3384 9580
rect 3332 9537 3341 9571
rect 3341 9537 3375 9571
rect 3375 9537 3384 9571
rect 3332 9528 3384 9537
rect 3700 9528 3752 9580
rect 5816 9596 5868 9648
rect 3884 9460 3936 9512
rect 3516 9392 3568 9444
rect 4160 9460 4212 9512
rect 4344 9503 4396 9512
rect 4344 9469 4353 9503
rect 4353 9469 4387 9503
rect 4387 9469 4396 9503
rect 4344 9460 4396 9469
rect 4436 9503 4488 9512
rect 4436 9469 4445 9503
rect 4445 9469 4479 9503
rect 4479 9469 4488 9503
rect 4436 9460 4488 9469
rect 5816 9460 5868 9512
rect 6460 9571 6512 9580
rect 6460 9537 6469 9571
rect 6469 9537 6503 9571
rect 6503 9537 6512 9571
rect 6460 9528 6512 9537
rect 6368 9460 6420 9512
rect 6920 9460 6972 9512
rect 7380 9528 7432 9580
rect 7564 9571 7616 9580
rect 7564 9537 7598 9571
rect 7598 9537 7616 9571
rect 7564 9528 7616 9537
rect 5172 9392 5224 9444
rect 2688 9324 2740 9376
rect 3240 9324 3292 9376
rect 3424 9324 3476 9376
rect 6276 9324 6328 9376
rect 7104 9324 7156 9376
rect 8392 9324 8444 9376
rect 1939 9222 1991 9274
rect 2003 9222 2055 9274
rect 2067 9222 2119 9274
rect 2131 9222 2183 9274
rect 2195 9222 2247 9274
rect 3917 9222 3969 9274
rect 3981 9222 4033 9274
rect 4045 9222 4097 9274
rect 4109 9222 4161 9274
rect 4173 9222 4225 9274
rect 5895 9222 5947 9274
rect 5959 9222 6011 9274
rect 6023 9222 6075 9274
rect 6087 9222 6139 9274
rect 6151 9222 6203 9274
rect 7873 9222 7925 9274
rect 7937 9222 7989 9274
rect 8001 9222 8053 9274
rect 8065 9222 8117 9274
rect 8129 9222 8181 9274
rect 2504 9120 2556 9172
rect 3332 9120 3384 9172
rect 5816 9163 5868 9172
rect 5816 9129 5825 9163
rect 5825 9129 5859 9163
rect 5859 9129 5868 9163
rect 5816 9120 5868 9129
rect 3148 8959 3200 8968
rect 3148 8925 3157 8959
rect 3157 8925 3191 8959
rect 3191 8925 3200 8959
rect 3148 8916 3200 8925
rect 3240 8959 3292 8968
rect 3240 8925 3249 8959
rect 3249 8925 3283 8959
rect 3283 8925 3292 8959
rect 3240 8916 3292 8925
rect 3516 8916 3568 8968
rect 4068 8916 4120 8968
rect 1676 8780 1728 8832
rect 4344 8848 4396 8900
rect 5724 8848 5776 8900
rect 7380 8959 7432 8968
rect 7380 8925 7389 8959
rect 7389 8925 7423 8959
rect 7423 8925 7432 8959
rect 7380 8916 7432 8925
rect 7656 8959 7708 8968
rect 7656 8925 7665 8959
rect 7665 8925 7699 8959
rect 7699 8925 7708 8959
rect 7656 8916 7708 8925
rect 8300 8916 8352 8968
rect 4252 8780 4304 8832
rect 5264 8780 5316 8832
rect 7748 8780 7800 8832
rect 2599 8678 2651 8730
rect 2663 8678 2715 8730
rect 2727 8678 2779 8730
rect 2791 8678 2843 8730
rect 2855 8678 2907 8730
rect 4577 8678 4629 8730
rect 4641 8678 4693 8730
rect 4705 8678 4757 8730
rect 4769 8678 4821 8730
rect 4833 8678 4885 8730
rect 6555 8678 6607 8730
rect 6619 8678 6671 8730
rect 6683 8678 6735 8730
rect 6747 8678 6799 8730
rect 6811 8678 6863 8730
rect 8533 8678 8585 8730
rect 8597 8678 8649 8730
rect 8661 8678 8713 8730
rect 8725 8678 8777 8730
rect 8789 8678 8841 8730
rect 2228 8576 2280 8628
rect 3148 8576 3200 8628
rect 3056 8508 3108 8560
rect 3332 8576 3384 8628
rect 5356 8576 5408 8628
rect 5816 8576 5868 8628
rect 7656 8576 7708 8628
rect 5080 8508 5132 8560
rect 1676 8483 1728 8492
rect 1676 8449 1685 8483
rect 1685 8449 1719 8483
rect 1719 8449 1728 8483
rect 1676 8440 1728 8449
rect 2320 8440 2372 8492
rect 2596 8440 2648 8492
rect 2872 8440 2924 8492
rect 3148 8440 3200 8492
rect 3240 8483 3292 8492
rect 3240 8449 3249 8483
rect 3249 8449 3283 8483
rect 3283 8449 3292 8483
rect 3240 8440 3292 8449
rect 3332 8483 3384 8492
rect 3332 8449 3341 8483
rect 3341 8449 3375 8483
rect 3375 8449 3384 8483
rect 3332 8440 3384 8449
rect 3424 8440 3476 8492
rect 4068 8440 4120 8492
rect 6736 8508 6788 8560
rect 5632 8440 5684 8492
rect 6644 8440 6696 8492
rect 7564 8483 7616 8492
rect 7564 8449 7598 8483
rect 7598 8449 7616 8483
rect 7564 8440 7616 8449
rect 5540 8415 5592 8424
rect 5540 8381 5549 8415
rect 5549 8381 5583 8415
rect 5583 8381 5592 8415
rect 5540 8372 5592 8381
rect 7288 8415 7340 8424
rect 7288 8381 7297 8415
rect 7297 8381 7331 8415
rect 7331 8381 7340 8415
rect 7288 8372 7340 8381
rect 5816 8304 5868 8356
rect 1584 8236 1636 8288
rect 2228 8236 2280 8288
rect 2596 8236 2648 8288
rect 3700 8236 3752 8288
rect 4436 8236 4488 8288
rect 5264 8236 5316 8288
rect 5448 8236 5500 8288
rect 6552 8304 6604 8356
rect 6368 8279 6420 8288
rect 6368 8245 6377 8279
rect 6377 8245 6411 8279
rect 6411 8245 6420 8279
rect 6368 8236 6420 8245
rect 7196 8236 7248 8288
rect 8392 8236 8444 8288
rect 8668 8279 8720 8288
rect 8668 8245 8677 8279
rect 8677 8245 8711 8279
rect 8711 8245 8720 8279
rect 8668 8236 8720 8245
rect 1939 8134 1991 8186
rect 2003 8134 2055 8186
rect 2067 8134 2119 8186
rect 2131 8134 2183 8186
rect 2195 8134 2247 8186
rect 3917 8134 3969 8186
rect 3981 8134 4033 8186
rect 4045 8134 4097 8186
rect 4109 8134 4161 8186
rect 4173 8134 4225 8186
rect 5895 8134 5947 8186
rect 5959 8134 6011 8186
rect 6023 8134 6075 8186
rect 6087 8134 6139 8186
rect 6151 8134 6203 8186
rect 7873 8134 7925 8186
rect 7937 8134 7989 8186
rect 8001 8134 8053 8186
rect 8065 8134 8117 8186
rect 8129 8134 8181 8186
rect 2872 7964 2924 8016
rect 3332 7896 3384 7948
rect 3700 7896 3752 7948
rect 5724 8075 5776 8084
rect 5724 8041 5733 8075
rect 5733 8041 5767 8075
rect 5767 8041 5776 8075
rect 5724 8032 5776 8041
rect 6368 8032 6420 8084
rect 6736 8032 6788 8084
rect 7196 8032 7248 8084
rect 7564 8032 7616 8084
rect 3884 7964 3936 8016
rect 5540 7964 5592 8016
rect 4988 7896 5040 7948
rect 5356 7896 5408 7948
rect 6184 7964 6236 8016
rect 2504 7803 2556 7812
rect 2504 7769 2522 7803
rect 2522 7769 2556 7803
rect 2504 7760 2556 7769
rect 2044 7692 2096 7744
rect 2412 7692 2464 7744
rect 4436 7828 4488 7880
rect 5080 7828 5132 7880
rect 6552 7896 6604 7948
rect 7380 7964 7432 8016
rect 7656 8007 7708 8016
rect 7656 7973 7665 8007
rect 7665 7973 7699 8007
rect 7699 7973 7708 8007
rect 7656 7964 7708 7973
rect 7748 7964 7800 8016
rect 6000 7803 6052 7812
rect 6000 7769 6009 7803
rect 6009 7769 6043 7803
rect 6043 7769 6052 7803
rect 6000 7760 6052 7769
rect 6092 7803 6144 7812
rect 6092 7769 6102 7803
rect 6102 7769 6136 7803
rect 6136 7769 6144 7803
rect 6092 7760 6144 7769
rect 6184 7760 6236 7812
rect 6644 7871 6696 7880
rect 6644 7837 6653 7871
rect 6653 7837 6687 7871
rect 6687 7837 6696 7871
rect 6644 7828 6696 7837
rect 7564 7896 7616 7948
rect 2964 7692 3016 7744
rect 3148 7692 3200 7744
rect 3424 7692 3476 7744
rect 3700 7692 3752 7744
rect 3792 7735 3844 7744
rect 3792 7701 3801 7735
rect 3801 7701 3835 7735
rect 3835 7701 3844 7735
rect 3792 7692 3844 7701
rect 4436 7735 4488 7744
rect 4436 7701 4445 7735
rect 4445 7701 4479 7735
rect 4479 7701 4488 7735
rect 4436 7692 4488 7701
rect 5080 7692 5132 7744
rect 6368 7692 6420 7744
rect 7012 7735 7064 7744
rect 7012 7701 7021 7735
rect 7021 7701 7055 7735
rect 7055 7701 7064 7735
rect 7012 7692 7064 7701
rect 7472 7803 7524 7812
rect 7472 7769 7481 7803
rect 7481 7769 7515 7803
rect 7515 7769 7524 7803
rect 7472 7760 7524 7769
rect 7564 7760 7616 7812
rect 8024 7828 8076 7880
rect 8392 7828 8444 7880
rect 8300 7760 8352 7812
rect 8116 7692 8168 7744
rect 8668 7692 8720 7744
rect 2599 7590 2651 7642
rect 2663 7590 2715 7642
rect 2727 7590 2779 7642
rect 2791 7590 2843 7642
rect 2855 7590 2907 7642
rect 4577 7590 4629 7642
rect 4641 7590 4693 7642
rect 4705 7590 4757 7642
rect 4769 7590 4821 7642
rect 4833 7590 4885 7642
rect 6555 7590 6607 7642
rect 6619 7590 6671 7642
rect 6683 7590 6735 7642
rect 6747 7590 6799 7642
rect 6811 7590 6863 7642
rect 8533 7590 8585 7642
rect 8597 7590 8649 7642
rect 8661 7590 8713 7642
rect 8725 7590 8777 7642
rect 8789 7590 8841 7642
rect 2412 7488 2464 7540
rect 2780 7488 2832 7540
rect 3332 7488 3384 7540
rect 3516 7488 3568 7540
rect 4344 7488 4396 7540
rect 7196 7488 7248 7540
rect 2044 7352 2096 7404
rect 3240 7352 3292 7404
rect 3792 7352 3844 7404
rect 1400 7191 1452 7200
rect 1400 7157 1409 7191
rect 1409 7157 1443 7191
rect 1443 7157 1452 7191
rect 1400 7148 1452 7157
rect 1584 7148 1636 7200
rect 2412 7284 2464 7336
rect 5264 7420 5316 7472
rect 4344 7395 4396 7404
rect 4344 7361 4353 7395
rect 4353 7361 4387 7395
rect 4387 7361 4396 7395
rect 4344 7352 4396 7361
rect 4620 7395 4672 7404
rect 4620 7361 4629 7395
rect 4629 7361 4663 7395
rect 4663 7361 4672 7395
rect 4620 7352 4672 7361
rect 4252 7284 4304 7336
rect 4528 7284 4580 7336
rect 4896 7352 4948 7404
rect 5908 7352 5960 7404
rect 5264 7284 5316 7336
rect 5448 7284 5500 7336
rect 5540 7284 5592 7336
rect 7104 7420 7156 7472
rect 7472 7420 7524 7472
rect 7840 7488 7892 7540
rect 8300 7488 8352 7540
rect 8208 7420 8260 7472
rect 6368 7352 6420 7404
rect 6828 7395 6880 7404
rect 6828 7361 6837 7395
rect 6837 7361 6871 7395
rect 6871 7361 6880 7395
rect 6828 7352 6880 7361
rect 6736 7327 6788 7336
rect 6736 7293 6745 7327
rect 6745 7293 6779 7327
rect 6779 7293 6788 7327
rect 6736 7284 6788 7293
rect 3240 7148 3292 7200
rect 4252 7148 4304 7200
rect 5172 7148 5224 7200
rect 6276 7148 6328 7200
rect 7840 7216 7892 7268
rect 7748 7191 7800 7200
rect 7748 7157 7757 7191
rect 7757 7157 7791 7191
rect 7791 7157 7800 7191
rect 7748 7148 7800 7157
rect 8300 7395 8352 7404
rect 8300 7361 8309 7395
rect 8309 7361 8343 7395
rect 8343 7361 8352 7395
rect 8300 7352 8352 7361
rect 8392 7216 8444 7268
rect 8484 7148 8536 7200
rect 1939 7046 1991 7098
rect 2003 7046 2055 7098
rect 2067 7046 2119 7098
rect 2131 7046 2183 7098
rect 2195 7046 2247 7098
rect 3917 7046 3969 7098
rect 3981 7046 4033 7098
rect 4045 7046 4097 7098
rect 4109 7046 4161 7098
rect 4173 7046 4225 7098
rect 5895 7046 5947 7098
rect 5959 7046 6011 7098
rect 6023 7046 6075 7098
rect 6087 7046 6139 7098
rect 6151 7046 6203 7098
rect 7873 7046 7925 7098
rect 7937 7046 7989 7098
rect 8001 7046 8053 7098
rect 8065 7046 8117 7098
rect 8129 7046 8181 7098
rect 6368 6944 6420 6996
rect 6736 6944 6788 6996
rect 8392 6944 8444 6996
rect 2780 6740 2832 6792
rect 1676 6715 1728 6724
rect 1676 6681 1710 6715
rect 1710 6681 1728 6715
rect 1676 6672 1728 6681
rect 3240 6876 3292 6928
rect 3884 6876 3936 6928
rect 4528 6876 4580 6928
rect 5540 6876 5592 6928
rect 5724 6876 5776 6928
rect 5816 6876 5868 6928
rect 6460 6876 6512 6928
rect 4896 6808 4948 6860
rect 3148 6740 3200 6792
rect 3516 6672 3568 6724
rect 3976 6783 4028 6792
rect 3976 6749 3985 6783
rect 3985 6749 4019 6783
rect 4019 6749 4028 6783
rect 3976 6740 4028 6749
rect 4068 6783 4120 6792
rect 4068 6749 4077 6783
rect 4077 6749 4111 6783
rect 4111 6749 4120 6783
rect 4068 6740 4120 6749
rect 4528 6783 4580 6792
rect 4528 6749 4537 6783
rect 4537 6749 4571 6783
rect 4571 6749 4580 6783
rect 4528 6740 4580 6749
rect 4620 6783 4672 6792
rect 4620 6749 4629 6783
rect 4629 6749 4663 6783
rect 4663 6749 4672 6783
rect 4620 6740 4672 6749
rect 1860 6604 1912 6656
rect 4068 6604 4120 6656
rect 5724 6783 5776 6792
rect 5724 6749 5733 6783
rect 5733 6749 5767 6783
rect 5767 6749 5776 6783
rect 5724 6740 5776 6749
rect 6184 6783 6236 6792
rect 6184 6749 6193 6783
rect 6193 6749 6227 6783
rect 6227 6749 6236 6783
rect 6184 6740 6236 6749
rect 6460 6783 6512 6792
rect 6460 6749 6469 6783
rect 6469 6749 6503 6783
rect 6503 6749 6512 6783
rect 6460 6740 6512 6749
rect 6920 6783 6972 6792
rect 6920 6749 6929 6783
rect 6929 6749 6963 6783
rect 6963 6749 6972 6783
rect 6920 6740 6972 6749
rect 7012 6740 7064 6792
rect 7472 6808 7524 6860
rect 8300 6808 8352 6860
rect 8944 6808 8996 6860
rect 7380 6740 7432 6792
rect 8208 6740 8260 6792
rect 9036 6740 9088 6792
rect 8116 6672 8168 6724
rect 5172 6604 5224 6656
rect 5448 6647 5500 6656
rect 5448 6613 5457 6647
rect 5457 6613 5491 6647
rect 5491 6613 5500 6647
rect 5448 6604 5500 6613
rect 6460 6604 6512 6656
rect 7012 6604 7064 6656
rect 7472 6647 7524 6656
rect 7472 6613 7481 6647
rect 7481 6613 7515 6647
rect 7515 6613 7524 6647
rect 7472 6604 7524 6613
rect 7656 6604 7708 6656
rect 7748 6604 7800 6656
rect 8392 6604 8444 6656
rect 2599 6502 2651 6554
rect 2663 6502 2715 6554
rect 2727 6502 2779 6554
rect 2791 6502 2843 6554
rect 2855 6502 2907 6554
rect 4577 6502 4629 6554
rect 4641 6502 4693 6554
rect 4705 6502 4757 6554
rect 4769 6502 4821 6554
rect 4833 6502 4885 6554
rect 6555 6502 6607 6554
rect 6619 6502 6671 6554
rect 6683 6502 6735 6554
rect 6747 6502 6799 6554
rect 6811 6502 6863 6554
rect 8533 6502 8585 6554
rect 8597 6502 8649 6554
rect 8661 6502 8713 6554
rect 8725 6502 8777 6554
rect 8789 6502 8841 6554
rect 1400 6332 1452 6384
rect 2412 6400 2464 6452
rect 2504 6443 2556 6452
rect 2504 6409 2513 6443
rect 2513 6409 2547 6443
rect 2547 6409 2556 6443
rect 2504 6400 2556 6409
rect 3332 6400 3384 6452
rect 1768 6264 1820 6316
rect 2320 6307 2372 6316
rect 2320 6273 2329 6307
rect 2329 6273 2363 6307
rect 2363 6273 2372 6307
rect 2320 6264 2372 6273
rect 2964 6332 3016 6384
rect 3608 6332 3660 6384
rect 3056 6264 3108 6316
rect 3516 6307 3568 6316
rect 3516 6273 3525 6307
rect 3525 6273 3559 6307
rect 3559 6273 3568 6307
rect 3516 6264 3568 6273
rect 3884 6264 3936 6316
rect 3976 6307 4028 6316
rect 3976 6273 3985 6307
rect 3985 6273 4019 6307
rect 4019 6273 4028 6307
rect 3976 6264 4028 6273
rect 1400 6103 1452 6112
rect 1400 6069 1409 6103
rect 1409 6069 1443 6103
rect 1443 6069 1452 6103
rect 1400 6060 1452 6069
rect 1768 6103 1820 6112
rect 1768 6069 1777 6103
rect 1777 6069 1811 6103
rect 1811 6069 1820 6103
rect 1768 6060 1820 6069
rect 4712 6400 4764 6452
rect 7380 6400 7432 6452
rect 7472 6400 7524 6452
rect 5632 6332 5684 6384
rect 5816 6332 5868 6384
rect 6184 6332 6236 6384
rect 4528 6264 4580 6316
rect 5724 6264 5776 6316
rect 6368 6307 6420 6316
rect 6368 6273 6377 6307
rect 6377 6273 6411 6307
rect 6411 6273 6420 6307
rect 6368 6264 6420 6273
rect 6920 6307 6972 6316
rect 6920 6273 6929 6307
rect 6929 6273 6963 6307
rect 6963 6273 6972 6307
rect 6920 6264 6972 6273
rect 7288 6307 7340 6316
rect 7288 6273 7297 6307
rect 7297 6273 7331 6307
rect 7331 6273 7340 6307
rect 7288 6264 7340 6273
rect 2228 6128 2280 6180
rect 3332 6060 3384 6112
rect 3608 6060 3660 6112
rect 4068 6060 4120 6112
rect 4344 6060 4396 6112
rect 6460 6060 6512 6112
rect 7288 6060 7340 6112
rect 7932 6060 7984 6112
rect 8944 6060 8996 6112
rect 1939 5958 1991 6010
rect 2003 5958 2055 6010
rect 2067 5958 2119 6010
rect 2131 5958 2183 6010
rect 2195 5958 2247 6010
rect 3917 5958 3969 6010
rect 3981 5958 4033 6010
rect 4045 5958 4097 6010
rect 4109 5958 4161 6010
rect 4173 5958 4225 6010
rect 5895 5958 5947 6010
rect 5959 5958 6011 6010
rect 6023 5958 6075 6010
rect 6087 5958 6139 6010
rect 6151 5958 6203 6010
rect 7873 5958 7925 6010
rect 7937 5958 7989 6010
rect 8001 5958 8053 6010
rect 8065 5958 8117 6010
rect 8129 5958 8181 6010
rect 1400 5856 1452 5908
rect 1676 5856 1728 5908
rect 1768 5856 1820 5908
rect 4620 5856 4672 5908
rect 5540 5856 5592 5908
rect 6000 5856 6052 5908
rect 7012 5899 7064 5908
rect 7012 5865 7021 5899
rect 7021 5865 7055 5899
rect 7055 5865 7064 5899
rect 7012 5856 7064 5865
rect 7564 5856 7616 5908
rect 7748 5856 7800 5908
rect 8208 5856 8260 5908
rect 3700 5720 3752 5772
rect 1860 5652 1912 5704
rect 2228 5652 2280 5704
rect 2320 5652 2372 5704
rect 2504 5652 2556 5704
rect 2872 5652 2924 5704
rect 3516 5652 3568 5704
rect 3240 5584 3292 5636
rect 3976 5652 4028 5704
rect 4068 5695 4120 5704
rect 4068 5661 4077 5695
rect 4077 5661 4111 5695
rect 4111 5661 4120 5695
rect 4068 5652 4120 5661
rect 4160 5652 4212 5704
rect 4252 5695 4304 5704
rect 4252 5661 4261 5695
rect 4261 5661 4295 5695
rect 4295 5661 4304 5695
rect 4252 5652 4304 5661
rect 4804 5720 4856 5772
rect 4712 5652 4764 5704
rect 4988 5652 5040 5704
rect 5172 5695 5224 5704
rect 5172 5661 5181 5695
rect 5181 5661 5215 5695
rect 5215 5661 5224 5695
rect 5172 5652 5224 5661
rect 5448 5720 5500 5772
rect 5816 5788 5868 5840
rect 5632 5720 5684 5772
rect 6460 5788 6512 5840
rect 8392 5788 8444 5840
rect 6460 5652 6512 5704
rect 6920 5695 6972 5704
rect 6920 5661 6929 5695
rect 6929 5661 6963 5695
rect 6963 5661 6972 5695
rect 6920 5652 6972 5661
rect 7012 5652 7064 5704
rect 7196 5652 7248 5704
rect 7656 5695 7708 5704
rect 7656 5661 7665 5695
rect 7665 5661 7699 5695
rect 7699 5661 7708 5695
rect 7656 5652 7708 5661
rect 8208 5652 8260 5704
rect 8392 5652 8444 5704
rect 1584 5516 1636 5568
rect 2504 5516 2556 5568
rect 2964 5516 3016 5568
rect 4160 5516 4212 5568
rect 4804 5516 4856 5568
rect 5356 5559 5408 5568
rect 5356 5525 5365 5559
rect 5365 5525 5399 5559
rect 5399 5525 5408 5559
rect 5356 5516 5408 5525
rect 5632 5516 5684 5568
rect 6276 5516 6328 5568
rect 7472 5559 7524 5568
rect 7472 5525 7481 5559
rect 7481 5525 7515 5559
rect 7515 5525 7524 5559
rect 7472 5516 7524 5525
rect 2599 5414 2651 5466
rect 2663 5414 2715 5466
rect 2727 5414 2779 5466
rect 2791 5414 2843 5466
rect 2855 5414 2907 5466
rect 4577 5414 4629 5466
rect 4641 5414 4693 5466
rect 4705 5414 4757 5466
rect 4769 5414 4821 5466
rect 4833 5414 4885 5466
rect 6555 5414 6607 5466
rect 6619 5414 6671 5466
rect 6683 5414 6735 5466
rect 6747 5414 6799 5466
rect 6811 5414 6863 5466
rect 8533 5414 8585 5466
rect 8597 5414 8649 5466
rect 8661 5414 8713 5466
rect 8725 5414 8777 5466
rect 8789 5414 8841 5466
rect 2872 5312 2924 5364
rect 4068 5312 4120 5364
rect 3056 5244 3108 5296
rect 3240 5287 3292 5296
rect 3240 5253 3249 5287
rect 3249 5253 3283 5287
rect 3283 5253 3292 5287
rect 3240 5244 3292 5253
rect 1400 5151 1452 5160
rect 1400 5117 1409 5151
rect 1409 5117 1443 5151
rect 1443 5117 1452 5151
rect 1400 5108 1452 5117
rect 2964 5176 3016 5228
rect 3700 5219 3752 5228
rect 3700 5185 3709 5219
rect 3709 5185 3743 5219
rect 3743 5185 3752 5219
rect 4620 5312 4672 5364
rect 4712 5312 4764 5364
rect 4252 5244 4304 5296
rect 5356 5312 5408 5364
rect 6368 5312 6420 5364
rect 6920 5312 6972 5364
rect 7472 5312 7524 5364
rect 3700 5176 3752 5185
rect 4436 5176 4488 5228
rect 5448 5244 5500 5296
rect 5724 5244 5776 5296
rect 3884 5108 3936 5160
rect 4252 5108 4304 5160
rect 4804 5176 4856 5228
rect 5356 5176 5408 5228
rect 5632 5219 5684 5228
rect 5632 5185 5641 5219
rect 5641 5185 5675 5219
rect 5675 5185 5684 5219
rect 5632 5176 5684 5185
rect 7564 5244 7616 5296
rect 8300 5244 8352 5296
rect 4160 5040 4212 5092
rect 1768 4972 1820 5024
rect 2596 4972 2648 5024
rect 3976 4972 4028 5024
rect 6184 5176 6236 5228
rect 6644 5176 6696 5228
rect 8208 5176 8260 5228
rect 8392 5219 8444 5228
rect 8392 5185 8401 5219
rect 8401 5185 8435 5219
rect 8435 5185 8444 5219
rect 8392 5176 8444 5185
rect 4988 5083 5040 5092
rect 4988 5049 4997 5083
rect 4997 5049 5031 5083
rect 5031 5049 5040 5083
rect 4988 5040 5040 5049
rect 5080 5040 5132 5092
rect 5816 5040 5868 5092
rect 7656 5108 7708 5160
rect 7748 5108 7800 5160
rect 5356 5015 5408 5024
rect 5356 4981 5365 5015
rect 5365 4981 5399 5015
rect 5399 4981 5408 5015
rect 5356 4972 5408 4981
rect 5448 4972 5500 5024
rect 6644 5083 6696 5092
rect 6644 5049 6653 5083
rect 6653 5049 6687 5083
rect 6687 5049 6696 5083
rect 6644 5040 6696 5049
rect 6000 4972 6052 5024
rect 6736 4972 6788 5024
rect 7564 5015 7616 5024
rect 7564 4981 7573 5015
rect 7573 4981 7607 5015
rect 7607 4981 7616 5015
rect 7564 4972 7616 4981
rect 1939 4870 1991 4922
rect 2003 4870 2055 4922
rect 2067 4870 2119 4922
rect 2131 4870 2183 4922
rect 2195 4870 2247 4922
rect 3917 4870 3969 4922
rect 3981 4870 4033 4922
rect 4045 4870 4097 4922
rect 4109 4870 4161 4922
rect 4173 4870 4225 4922
rect 5895 4870 5947 4922
rect 5959 4870 6011 4922
rect 6023 4870 6075 4922
rect 6087 4870 6139 4922
rect 6151 4870 6203 4922
rect 7873 4870 7925 4922
rect 7937 4870 7989 4922
rect 8001 4870 8053 4922
rect 8065 4870 8117 4922
rect 8129 4870 8181 4922
rect 1768 4768 1820 4820
rect 3056 4768 3108 4820
rect 3148 4768 3200 4820
rect 2320 4675 2372 4684
rect 2320 4641 2329 4675
rect 2329 4641 2363 4675
rect 2363 4641 2372 4675
rect 2320 4632 2372 4641
rect 3516 4700 3568 4752
rect 3976 4768 4028 4820
rect 5172 4811 5224 4820
rect 5172 4777 5181 4811
rect 5181 4777 5215 4811
rect 5215 4777 5224 4811
rect 5172 4768 5224 4777
rect 5448 4700 5500 4752
rect 6460 4811 6512 4820
rect 6460 4777 6469 4811
rect 6469 4777 6503 4811
rect 6503 4777 6512 4811
rect 6460 4768 6512 4777
rect 6736 4811 6788 4820
rect 6736 4777 6745 4811
rect 6745 4777 6779 4811
rect 6779 4777 6788 4811
rect 6736 4768 6788 4777
rect 7012 4768 7064 4820
rect 7472 4768 7524 4820
rect 8208 4768 8260 4820
rect 4436 4632 4488 4684
rect 1952 4539 2004 4548
rect 1952 4505 1961 4539
rect 1961 4505 1995 4539
rect 1995 4505 2004 4539
rect 1952 4496 2004 4505
rect 3056 4564 3108 4616
rect 2136 4471 2188 4480
rect 2136 4437 2145 4471
rect 2145 4437 2179 4471
rect 2179 4437 2188 4471
rect 2136 4428 2188 4437
rect 2596 4471 2648 4480
rect 2596 4437 2605 4471
rect 2605 4437 2639 4471
rect 2639 4437 2648 4471
rect 2596 4428 2648 4437
rect 2872 4496 2924 4548
rect 3424 4564 3476 4616
rect 4068 4607 4120 4616
rect 4068 4573 4077 4607
rect 4077 4573 4111 4607
rect 4111 4573 4120 4607
rect 4068 4564 4120 4573
rect 3240 4428 3292 4480
rect 3332 4471 3384 4480
rect 3332 4437 3341 4471
rect 3341 4437 3375 4471
rect 3375 4437 3384 4471
rect 3332 4428 3384 4437
rect 4068 4428 4120 4480
rect 4252 4471 4304 4480
rect 4252 4437 4261 4471
rect 4261 4437 4295 4471
rect 4295 4437 4304 4471
rect 4252 4428 4304 4437
rect 4528 4607 4580 4616
rect 4528 4573 4537 4607
rect 4537 4573 4571 4607
rect 4571 4573 4580 4607
rect 4528 4564 4580 4573
rect 5080 4632 5132 4684
rect 5632 4607 5684 4616
rect 5632 4573 5641 4607
rect 5641 4573 5675 4607
rect 5675 4573 5684 4607
rect 5632 4564 5684 4573
rect 4896 4496 4948 4548
rect 4528 4428 4580 4480
rect 4712 4428 4764 4480
rect 5448 4496 5500 4548
rect 5540 4428 5592 4480
rect 6184 4632 6236 4684
rect 6460 4607 6512 4616
rect 6460 4573 6469 4607
rect 6469 4573 6503 4607
rect 6503 4573 6512 4607
rect 6460 4564 6512 4573
rect 7012 4607 7064 4616
rect 7012 4573 7021 4607
rect 7021 4573 7055 4607
rect 7055 4573 7064 4607
rect 7012 4564 7064 4573
rect 7196 4607 7248 4616
rect 7196 4573 7205 4607
rect 7205 4573 7239 4607
rect 7239 4573 7248 4607
rect 7196 4564 7248 4573
rect 8300 4607 8352 4616
rect 8300 4573 8309 4607
rect 8309 4573 8343 4607
rect 8343 4573 8352 4607
rect 8300 4564 8352 4573
rect 5908 4471 5960 4480
rect 5908 4437 5917 4471
rect 5917 4437 5951 4471
rect 5951 4437 5960 4471
rect 5908 4428 5960 4437
rect 6000 4471 6052 4480
rect 6000 4437 6009 4471
rect 6009 4437 6043 4471
rect 6043 4437 6052 4471
rect 6000 4428 6052 4437
rect 6184 4428 6236 4480
rect 6828 4471 6880 4480
rect 6828 4437 6837 4471
rect 6837 4437 6871 4471
rect 6871 4437 6880 4471
rect 6828 4428 6880 4437
rect 7104 4539 7156 4548
rect 7104 4505 7113 4539
rect 7113 4505 7147 4539
rect 7147 4505 7156 4539
rect 7104 4496 7156 4505
rect 8576 4539 8628 4548
rect 8576 4505 8585 4539
rect 8585 4505 8619 4539
rect 8619 4505 8628 4539
rect 8576 4496 8628 4505
rect 2599 4326 2651 4378
rect 2663 4326 2715 4378
rect 2727 4326 2779 4378
rect 2791 4326 2843 4378
rect 2855 4326 2907 4378
rect 4577 4326 4629 4378
rect 4641 4326 4693 4378
rect 4705 4326 4757 4378
rect 4769 4326 4821 4378
rect 4833 4326 4885 4378
rect 6555 4326 6607 4378
rect 6619 4326 6671 4378
rect 6683 4326 6735 4378
rect 6747 4326 6799 4378
rect 6811 4326 6863 4378
rect 8533 4326 8585 4378
rect 8597 4326 8649 4378
rect 8661 4326 8713 4378
rect 8725 4326 8777 4378
rect 8789 4326 8841 4378
rect 1952 4224 2004 4276
rect 1492 4131 1544 4140
rect 1492 4097 1501 4131
rect 1501 4097 1535 4131
rect 1535 4097 1544 4131
rect 1492 4088 1544 4097
rect 1676 4131 1728 4140
rect 1676 4097 1685 4131
rect 1685 4097 1719 4131
rect 1719 4097 1728 4131
rect 1676 4088 1728 4097
rect 1768 3952 1820 4004
rect 1860 3927 1912 3936
rect 1860 3893 1869 3927
rect 1869 3893 1903 3927
rect 1903 3893 1912 3927
rect 1860 3884 1912 3893
rect 2228 4131 2280 4140
rect 2228 4097 2237 4131
rect 2237 4097 2271 4131
rect 2271 4097 2280 4131
rect 2228 4088 2280 4097
rect 2320 4020 2372 4072
rect 3976 4156 4028 4208
rect 2964 4088 3016 4140
rect 3792 4088 3844 4140
rect 4160 4224 4212 4276
rect 5908 4224 5960 4276
rect 7104 4224 7156 4276
rect 8392 4224 8444 4276
rect 4988 4131 5040 4140
rect 4988 4097 4997 4131
rect 4997 4097 5031 4131
rect 5031 4097 5040 4131
rect 4988 4088 5040 4097
rect 2872 3952 2924 4004
rect 3240 3952 3292 4004
rect 4528 4020 4580 4072
rect 4068 3952 4120 4004
rect 5540 4156 5592 4208
rect 5632 4088 5684 4140
rect 6276 4088 6328 4140
rect 6184 4020 6236 4072
rect 2412 3884 2464 3936
rect 2504 3927 2556 3936
rect 2504 3893 2513 3927
rect 2513 3893 2547 3927
rect 2547 3893 2556 3927
rect 2504 3884 2556 3893
rect 5540 3884 5592 3936
rect 5632 3927 5684 3936
rect 5632 3893 5641 3927
rect 5641 3893 5675 3927
rect 5675 3893 5684 3927
rect 5632 3884 5684 3893
rect 6368 3884 6420 3936
rect 6828 4088 6880 4140
rect 7104 4088 7156 4140
rect 7564 4088 7616 4140
rect 8944 4088 8996 4140
rect 8300 4020 8352 4072
rect 6736 3952 6788 4004
rect 7012 3952 7064 4004
rect 7196 3884 7248 3936
rect 1939 3782 1991 3834
rect 2003 3782 2055 3834
rect 2067 3782 2119 3834
rect 2131 3782 2183 3834
rect 2195 3782 2247 3834
rect 3917 3782 3969 3834
rect 3981 3782 4033 3834
rect 4045 3782 4097 3834
rect 4109 3782 4161 3834
rect 4173 3782 4225 3834
rect 5895 3782 5947 3834
rect 5959 3782 6011 3834
rect 6023 3782 6075 3834
rect 6087 3782 6139 3834
rect 6151 3782 6203 3834
rect 7873 3782 7925 3834
rect 7937 3782 7989 3834
rect 8001 3782 8053 3834
rect 8065 3782 8117 3834
rect 8129 3782 8181 3834
rect 2504 3680 2556 3732
rect 2872 3723 2924 3732
rect 2872 3689 2881 3723
rect 2881 3689 2915 3723
rect 2915 3689 2924 3723
rect 2872 3680 2924 3689
rect 1400 3587 1452 3596
rect 1400 3553 1409 3587
rect 1409 3553 1443 3587
rect 1443 3553 1452 3587
rect 1400 3544 1452 3553
rect 3424 3680 3476 3732
rect 3608 3680 3660 3732
rect 3700 3680 3752 3732
rect 4620 3680 4672 3732
rect 5540 3680 5592 3732
rect 7472 3680 7524 3732
rect 3332 3655 3384 3664
rect 3332 3621 3341 3655
rect 3341 3621 3375 3655
rect 3375 3621 3384 3655
rect 3332 3612 3384 3621
rect 2964 3544 3016 3596
rect 3056 3587 3108 3596
rect 3056 3553 3065 3587
rect 3065 3553 3099 3587
rect 3099 3553 3108 3587
rect 3056 3544 3108 3553
rect 5172 3655 5224 3664
rect 5172 3621 5181 3655
rect 5181 3621 5215 3655
rect 5215 3621 5224 3655
rect 5172 3612 5224 3621
rect 3240 3519 3292 3528
rect 3240 3485 3249 3519
rect 3249 3485 3283 3519
rect 3283 3485 3292 3519
rect 3240 3476 3292 3485
rect 3884 3476 3936 3528
rect 3424 3408 3476 3460
rect 3056 3340 3108 3392
rect 3792 3340 3844 3392
rect 3884 3383 3936 3392
rect 3884 3349 3893 3383
rect 3893 3349 3927 3383
rect 3927 3349 3936 3383
rect 3884 3340 3936 3349
rect 3976 3383 4028 3392
rect 3976 3349 3985 3383
rect 3985 3349 4019 3383
rect 4019 3349 4028 3383
rect 3976 3340 4028 3349
rect 4068 3383 4120 3392
rect 4068 3349 4077 3383
rect 4077 3349 4111 3383
rect 4111 3349 4120 3383
rect 4068 3340 4120 3349
rect 4436 3476 4488 3528
rect 4528 3519 4580 3528
rect 4528 3485 4537 3519
rect 4537 3485 4571 3519
rect 4571 3485 4580 3519
rect 4528 3476 4580 3485
rect 4620 3519 4672 3528
rect 4620 3485 4629 3519
rect 4629 3485 4663 3519
rect 4663 3485 4672 3519
rect 4620 3476 4672 3485
rect 4988 3476 5040 3528
rect 5172 3476 5224 3528
rect 5264 3476 5316 3528
rect 6736 3544 6788 3596
rect 4620 3340 4672 3392
rect 4988 3383 5040 3392
rect 4988 3349 4997 3383
rect 4997 3349 5031 3383
rect 5031 3349 5040 3383
rect 4988 3340 5040 3349
rect 6276 3408 6328 3460
rect 7104 3476 7156 3528
rect 7012 3340 7064 3392
rect 7288 3408 7340 3460
rect 2599 3238 2651 3290
rect 2663 3238 2715 3290
rect 2727 3238 2779 3290
rect 2791 3238 2843 3290
rect 2855 3238 2907 3290
rect 4577 3238 4629 3290
rect 4641 3238 4693 3290
rect 4705 3238 4757 3290
rect 4769 3238 4821 3290
rect 4833 3238 4885 3290
rect 6555 3238 6607 3290
rect 6619 3238 6671 3290
rect 6683 3238 6735 3290
rect 6747 3238 6799 3290
rect 6811 3238 6863 3290
rect 8533 3238 8585 3290
rect 8597 3238 8649 3290
rect 8661 3238 8713 3290
rect 8725 3238 8777 3290
rect 8789 3238 8841 3290
rect 1400 3136 1452 3188
rect 1860 3136 1912 3188
rect 2780 3068 2832 3120
rect 1768 3043 1820 3052
rect 1768 3009 1795 3043
rect 1795 3009 1820 3043
rect 1768 3000 1820 3009
rect 2044 3043 2096 3052
rect 2044 3009 2053 3043
rect 2053 3009 2087 3043
rect 2087 3009 2096 3043
rect 2044 3000 2096 3009
rect 3608 3000 3660 3052
rect 4160 3136 4212 3188
rect 4896 3136 4948 3188
rect 4988 3136 5040 3188
rect 4344 3111 4396 3120
rect 4344 3077 4353 3111
rect 4353 3077 4387 3111
rect 4387 3077 4396 3111
rect 4344 3068 4396 3077
rect 5632 3136 5684 3188
rect 6736 3136 6788 3188
rect 6920 3136 6972 3188
rect 7012 3136 7064 3188
rect 5540 3068 5592 3120
rect 3240 2864 3292 2916
rect 4988 2975 5040 2984
rect 4988 2941 4997 2975
rect 4997 2941 5031 2975
rect 5031 2941 5040 2975
rect 4988 2932 5040 2941
rect 5632 2975 5684 2984
rect 5632 2941 5641 2975
rect 5641 2941 5675 2975
rect 5675 2941 5684 2975
rect 5632 2932 5684 2941
rect 5908 3000 5960 3052
rect 7380 3068 7432 3120
rect 6920 3043 6972 3052
rect 6920 3009 6929 3043
rect 6929 3009 6963 3043
rect 6963 3009 6972 3043
rect 6920 3000 6972 3009
rect 7196 3043 7248 3052
rect 7196 3009 7205 3043
rect 7205 3009 7239 3043
rect 7239 3009 7248 3043
rect 7196 3000 7248 3009
rect 8024 3179 8076 3188
rect 8024 3145 8033 3179
rect 8033 3145 8067 3179
rect 8067 3145 8076 3179
rect 8024 3136 8076 3145
rect 7748 3000 7800 3052
rect 8300 3136 8352 3188
rect 5816 2864 5868 2916
rect 20 2796 72 2848
rect 2320 2796 2372 2848
rect 2596 2796 2648 2848
rect 5172 2839 5224 2848
rect 5172 2805 5181 2839
rect 5181 2805 5215 2839
rect 5215 2805 5224 2839
rect 5172 2796 5224 2805
rect 6368 2796 6420 2848
rect 7012 2864 7064 2916
rect 8484 2932 8536 2984
rect 6828 2796 6880 2848
rect 7656 2796 7708 2848
rect 8300 2796 8352 2848
rect 1939 2694 1991 2746
rect 2003 2694 2055 2746
rect 2067 2694 2119 2746
rect 2131 2694 2183 2746
rect 2195 2694 2247 2746
rect 3917 2694 3969 2746
rect 3981 2694 4033 2746
rect 4045 2694 4097 2746
rect 4109 2694 4161 2746
rect 4173 2694 4225 2746
rect 5895 2694 5947 2746
rect 5959 2694 6011 2746
rect 6023 2694 6075 2746
rect 6087 2694 6139 2746
rect 6151 2694 6203 2746
rect 7873 2694 7925 2746
rect 7937 2694 7989 2746
rect 8001 2694 8053 2746
rect 8065 2694 8117 2746
rect 8129 2694 8181 2746
rect 1768 2592 1820 2644
rect 2504 2592 2556 2644
rect 2780 2592 2832 2644
rect 3608 2592 3660 2644
rect 4988 2592 5040 2644
rect 5632 2592 5684 2644
rect 5908 2592 5960 2644
rect 6276 2592 6328 2644
rect 7012 2635 7064 2644
rect 7012 2601 7021 2635
rect 7021 2601 7055 2635
rect 7055 2601 7064 2635
rect 7012 2592 7064 2601
rect 3240 2456 3292 2508
rect 3332 2431 3384 2440
rect 3332 2397 3341 2431
rect 3341 2397 3375 2431
rect 3375 2397 3384 2431
rect 3332 2388 3384 2397
rect 3424 2431 3476 2440
rect 3424 2397 3433 2431
rect 3433 2397 3467 2431
rect 3467 2397 3476 2431
rect 3424 2388 3476 2397
rect 3056 2363 3108 2372
rect 3056 2329 3065 2363
rect 3065 2329 3099 2363
rect 3099 2329 3108 2363
rect 3056 2320 3108 2329
rect 3516 2295 3568 2304
rect 3516 2261 3525 2295
rect 3525 2261 3559 2295
rect 3559 2261 3568 2295
rect 3516 2252 3568 2261
rect 5264 2431 5316 2440
rect 5264 2397 5273 2431
rect 5273 2397 5307 2431
rect 5307 2397 5316 2431
rect 5264 2388 5316 2397
rect 5540 2431 5592 2440
rect 5540 2397 5549 2431
rect 5549 2397 5583 2431
rect 5583 2397 5592 2431
rect 5540 2388 5592 2397
rect 5632 2388 5684 2440
rect 6460 2524 6512 2576
rect 6828 2524 6880 2576
rect 6368 2499 6420 2508
rect 6368 2465 6377 2499
rect 6377 2465 6411 2499
rect 6411 2465 6420 2499
rect 6368 2456 6420 2465
rect 7656 2524 7708 2576
rect 5816 2431 5868 2440
rect 5816 2397 5825 2431
rect 5825 2397 5859 2431
rect 5859 2397 5868 2431
rect 5816 2388 5868 2397
rect 5908 2431 5960 2440
rect 5908 2397 5917 2431
rect 5917 2397 5951 2431
rect 5951 2397 5960 2431
rect 5908 2388 5960 2397
rect 6736 2431 6788 2440
rect 6736 2397 6745 2431
rect 6745 2397 6779 2431
rect 6779 2397 6788 2431
rect 6736 2388 6788 2397
rect 4252 2320 4304 2372
rect 5172 2320 5224 2372
rect 7196 2431 7248 2440
rect 7196 2397 7205 2431
rect 7205 2397 7239 2431
rect 7239 2397 7248 2431
rect 7196 2388 7248 2397
rect 7932 2431 7984 2440
rect 7932 2397 7941 2431
rect 7941 2397 7975 2431
rect 7975 2397 7984 2431
rect 7932 2388 7984 2397
rect 8300 2524 8352 2576
rect 8484 2524 8536 2576
rect 6460 2295 6512 2304
rect 6460 2261 6469 2295
rect 6469 2261 6503 2295
rect 6503 2261 6512 2295
rect 6460 2252 6512 2261
rect 7472 2295 7524 2304
rect 7472 2261 7481 2295
rect 7481 2261 7515 2295
rect 7515 2261 7524 2295
rect 7472 2252 7524 2261
rect 8024 2295 8076 2304
rect 8024 2261 8033 2295
rect 8033 2261 8067 2295
rect 8067 2261 8076 2295
rect 8024 2252 8076 2261
rect 2599 2150 2651 2202
rect 2663 2150 2715 2202
rect 2727 2150 2779 2202
rect 2791 2150 2843 2202
rect 2855 2150 2907 2202
rect 4577 2150 4629 2202
rect 4641 2150 4693 2202
rect 4705 2150 4757 2202
rect 4769 2150 4821 2202
rect 4833 2150 4885 2202
rect 6555 2150 6607 2202
rect 6619 2150 6671 2202
rect 6683 2150 6735 2202
rect 6747 2150 6799 2202
rect 6811 2150 6863 2202
rect 8533 2150 8585 2202
rect 8597 2150 8649 2202
rect 8661 2150 8713 2202
rect 8725 2150 8777 2202
rect 8789 2150 8841 2202
rect 1584 1844 1636 1896
rect 8024 2048 8076 2100
rect 3056 1980 3108 2032
rect 5356 1980 5408 2032
rect 5724 1980 5776 2032
rect 3516 1912 3568 1964
rect 3792 1844 3844 1896
rect 6460 1844 6512 1896
rect 3700 1708 3752 1760
rect 7472 1708 7524 1760
<< metal2 >>
rect 5814 11556 5870 12356
rect 2599 9820 2907 9829
rect 2599 9818 2605 9820
rect 2661 9818 2685 9820
rect 2741 9818 2765 9820
rect 2821 9818 2845 9820
rect 2901 9818 2907 9820
rect 2661 9766 2663 9818
rect 2843 9766 2845 9818
rect 2599 9764 2605 9766
rect 2661 9764 2685 9766
rect 2741 9764 2765 9766
rect 2821 9764 2845 9766
rect 2901 9764 2907 9766
rect 2599 9755 2907 9764
rect 4577 9820 4885 9829
rect 4577 9818 4583 9820
rect 4639 9818 4663 9820
rect 4719 9818 4743 9820
rect 4799 9818 4823 9820
rect 4879 9818 4885 9820
rect 4639 9766 4641 9818
rect 4821 9766 4823 9818
rect 4577 9764 4583 9766
rect 4639 9764 4663 9766
rect 4719 9764 4743 9766
rect 4799 9764 4823 9766
rect 4879 9764 4885 9766
rect 4577 9755 4885 9764
rect 2688 9716 2740 9722
rect 2688 9658 2740 9664
rect 2044 9648 2096 9654
rect 2044 9590 2096 9596
rect 2056 9518 2084 9590
rect 1676 9512 1728 9518
rect 1676 9454 1728 9460
rect 2044 9512 2096 9518
rect 2044 9454 2096 9460
rect 2320 9512 2372 9518
rect 2320 9454 2372 9460
rect 2412 9512 2464 9518
rect 2412 9454 2464 9460
rect 1688 8838 1716 9454
rect 1860 9376 1912 9382
rect 1860 9318 1912 9324
rect 1676 8832 1728 8838
rect 1676 8774 1728 8780
rect 1688 8498 1716 8774
rect 1676 8492 1728 8498
rect 1676 8434 1728 8440
rect 1584 8288 1636 8294
rect 1584 8230 1636 8236
rect 1596 7206 1624 8230
rect 1400 7200 1452 7206
rect 1400 7142 1452 7148
rect 1584 7200 1636 7206
rect 1584 7142 1636 7148
rect 1412 6390 1440 7142
rect 1400 6384 1452 6390
rect 1400 6326 1452 6332
rect 1400 6112 1452 6118
rect 1400 6054 1452 6060
rect 1412 5914 1440 6054
rect 1400 5908 1452 5914
rect 1400 5850 1452 5856
rect 1596 5574 1624 7142
rect 1872 6984 1900 9318
rect 1939 9276 2247 9285
rect 1939 9274 1945 9276
rect 2001 9274 2025 9276
rect 2081 9274 2105 9276
rect 2161 9274 2185 9276
rect 2241 9274 2247 9276
rect 2001 9222 2003 9274
rect 2183 9222 2185 9274
rect 1939 9220 1945 9222
rect 2001 9220 2025 9222
rect 2081 9220 2105 9222
rect 2161 9220 2185 9222
rect 2241 9220 2247 9222
rect 1939 9211 2247 9220
rect 2228 8628 2280 8634
rect 2228 8570 2280 8576
rect 2240 8294 2268 8570
rect 2332 8498 2360 9454
rect 2424 9160 2452 9454
rect 2700 9382 2728 9658
rect 5828 9654 5856 11556
rect 6555 9820 6863 9829
rect 6555 9818 6561 9820
rect 6617 9818 6641 9820
rect 6697 9818 6721 9820
rect 6777 9818 6801 9820
rect 6857 9818 6863 9820
rect 6617 9766 6619 9818
rect 6799 9766 6801 9818
rect 6555 9764 6561 9766
rect 6617 9764 6641 9766
rect 6697 9764 6721 9766
rect 6777 9764 6801 9766
rect 6857 9764 6863 9766
rect 6555 9755 6863 9764
rect 8533 9820 8841 9829
rect 8533 9818 8539 9820
rect 8595 9818 8619 9820
rect 8675 9818 8699 9820
rect 8755 9818 8779 9820
rect 8835 9818 8841 9820
rect 8595 9766 8597 9818
rect 8777 9766 8779 9818
rect 8533 9764 8539 9766
rect 8595 9764 8619 9766
rect 8675 9764 8699 9766
rect 8755 9764 8779 9766
rect 8835 9764 8841 9766
rect 8533 9755 8841 9764
rect 5816 9648 5868 9654
rect 5816 9590 5868 9596
rect 3332 9580 3384 9586
rect 3332 9522 3384 9528
rect 3700 9580 3752 9586
rect 3700 9522 3752 9528
rect 6460 9580 6512 9586
rect 6460 9522 6512 9528
rect 7380 9580 7432 9586
rect 7380 9522 7432 9528
rect 7564 9580 7616 9586
rect 7564 9522 7616 9528
rect 2688 9376 2740 9382
rect 2688 9318 2740 9324
rect 3240 9376 3292 9382
rect 3240 9318 3292 9324
rect 2504 9172 2556 9178
rect 2424 9132 2504 9160
rect 2504 9114 2556 9120
rect 3252 8974 3280 9318
rect 3344 9178 3372 9522
rect 3516 9444 3568 9450
rect 3516 9386 3568 9392
rect 3424 9376 3476 9382
rect 3424 9318 3476 9324
rect 3332 9172 3384 9178
rect 3332 9114 3384 9120
rect 3148 8968 3200 8974
rect 3148 8910 3200 8916
rect 3240 8968 3292 8974
rect 3240 8910 3292 8916
rect 2599 8732 2907 8741
rect 2599 8730 2605 8732
rect 2661 8730 2685 8732
rect 2741 8730 2765 8732
rect 2821 8730 2845 8732
rect 2901 8730 2907 8732
rect 2661 8678 2663 8730
rect 2843 8678 2845 8730
rect 2599 8676 2605 8678
rect 2661 8676 2685 8678
rect 2741 8676 2765 8678
rect 2821 8676 2845 8678
rect 2901 8676 2907 8678
rect 2599 8667 2907 8676
rect 3160 8634 3188 8910
rect 3344 8634 3372 9114
rect 3148 8628 3200 8634
rect 3148 8570 3200 8576
rect 3332 8628 3384 8634
rect 3332 8570 3384 8576
rect 3056 8560 3108 8566
rect 3056 8502 3108 8508
rect 2320 8492 2372 8498
rect 2320 8434 2372 8440
rect 2596 8492 2648 8498
rect 2596 8434 2648 8440
rect 2872 8492 2924 8498
rect 2872 8434 2924 8440
rect 2608 8294 2636 8434
rect 2228 8288 2280 8294
rect 2228 8230 2280 8236
rect 2596 8288 2648 8294
rect 2596 8230 2648 8236
rect 1939 8188 2247 8197
rect 1939 8186 1945 8188
rect 2001 8186 2025 8188
rect 2081 8186 2105 8188
rect 2161 8186 2185 8188
rect 2241 8186 2247 8188
rect 2001 8134 2003 8186
rect 2183 8134 2185 8186
rect 1939 8132 1945 8134
rect 2001 8132 2025 8134
rect 2081 8132 2105 8134
rect 2161 8132 2185 8134
rect 2241 8132 2247 8134
rect 1939 8123 2247 8132
rect 2884 8022 2912 8434
rect 2872 8016 2924 8022
rect 2872 7958 2924 7964
rect 2504 7812 2556 7818
rect 2504 7754 2556 7760
rect 2044 7744 2096 7750
rect 2044 7686 2096 7692
rect 2412 7744 2464 7750
rect 2412 7686 2464 7692
rect 2056 7410 2084 7686
rect 2424 7546 2452 7686
rect 2412 7540 2464 7546
rect 2412 7482 2464 7488
rect 2044 7404 2096 7410
rect 2044 7346 2096 7352
rect 2412 7336 2464 7342
rect 2412 7278 2464 7284
rect 1939 7100 2247 7109
rect 1939 7098 1945 7100
rect 2001 7098 2025 7100
rect 2081 7098 2105 7100
rect 2161 7098 2185 7100
rect 2241 7098 2247 7100
rect 2001 7046 2003 7098
rect 2183 7046 2185 7098
rect 1939 7044 1945 7046
rect 2001 7044 2025 7046
rect 2081 7044 2105 7046
rect 2161 7044 2185 7046
rect 2241 7044 2247 7046
rect 1939 7035 2247 7044
rect 1872 6956 2268 6984
rect 1676 6724 1728 6730
rect 1676 6666 1728 6672
rect 1688 5914 1716 6666
rect 1860 6656 1912 6662
rect 1860 6598 1912 6604
rect 1766 6352 1822 6361
rect 1766 6287 1768 6296
rect 1820 6287 1822 6296
rect 1768 6258 1820 6264
rect 1768 6112 1820 6118
rect 1768 6054 1820 6060
rect 1780 5914 1808 6054
rect 1676 5908 1728 5914
rect 1676 5850 1728 5856
rect 1768 5908 1820 5914
rect 1768 5850 1820 5856
rect 1872 5710 1900 6598
rect 2240 6186 2268 6956
rect 2424 6458 2452 7278
rect 2516 6458 2544 7754
rect 2964 7744 3016 7750
rect 2964 7686 3016 7692
rect 2599 7644 2907 7653
rect 2599 7642 2605 7644
rect 2661 7642 2685 7644
rect 2741 7642 2765 7644
rect 2821 7642 2845 7644
rect 2901 7642 2907 7644
rect 2661 7590 2663 7642
rect 2843 7590 2845 7642
rect 2599 7588 2605 7590
rect 2661 7588 2685 7590
rect 2741 7588 2765 7590
rect 2821 7588 2845 7590
rect 2901 7588 2907 7590
rect 2599 7579 2907 7588
rect 2780 7540 2832 7546
rect 2780 7482 2832 7488
rect 2792 6798 2820 7482
rect 2780 6792 2832 6798
rect 2780 6734 2832 6740
rect 2599 6556 2907 6565
rect 2599 6554 2605 6556
rect 2661 6554 2685 6556
rect 2741 6554 2765 6556
rect 2821 6554 2845 6556
rect 2901 6554 2907 6556
rect 2661 6502 2663 6554
rect 2843 6502 2845 6554
rect 2599 6500 2605 6502
rect 2661 6500 2685 6502
rect 2741 6500 2765 6502
rect 2821 6500 2845 6502
rect 2901 6500 2907 6502
rect 2599 6491 2907 6500
rect 2412 6452 2464 6458
rect 2412 6394 2464 6400
rect 2504 6452 2556 6458
rect 2504 6394 2556 6400
rect 2976 6390 3004 7686
rect 3068 6780 3096 8502
rect 3436 8498 3464 9318
rect 3528 8974 3556 9386
rect 3516 8968 3568 8974
rect 3516 8910 3568 8916
rect 3606 8936 3662 8945
rect 3606 8871 3662 8880
rect 3148 8492 3200 8498
rect 3148 8434 3200 8440
rect 3240 8492 3292 8498
rect 3240 8434 3292 8440
rect 3332 8492 3384 8498
rect 3332 8434 3384 8440
rect 3424 8492 3476 8498
rect 3424 8434 3476 8440
rect 3160 7750 3188 8434
rect 3148 7744 3200 7750
rect 3148 7686 3200 7692
rect 3252 7410 3280 8434
rect 3344 7954 3372 8434
rect 3332 7948 3384 7954
rect 3332 7890 3384 7896
rect 3344 7546 3372 7890
rect 3424 7744 3476 7750
rect 3424 7686 3476 7692
rect 3332 7540 3384 7546
rect 3332 7482 3384 7488
rect 3436 7426 3464 7686
rect 3516 7540 3568 7546
rect 3516 7482 3568 7488
rect 3240 7404 3292 7410
rect 3240 7346 3292 7352
rect 3344 7398 3464 7426
rect 3240 7200 3292 7206
rect 3240 7142 3292 7148
rect 3252 6934 3280 7142
rect 3240 6928 3292 6934
rect 3240 6870 3292 6876
rect 3148 6792 3200 6798
rect 3068 6752 3148 6780
rect 2964 6384 3016 6390
rect 2964 6326 3016 6332
rect 3068 6322 3096 6752
rect 3148 6734 3200 6740
rect 3344 6458 3372 7398
rect 3528 6848 3556 7482
rect 3436 6820 3556 6848
rect 3332 6452 3384 6458
rect 3332 6394 3384 6400
rect 2320 6316 2372 6322
rect 2320 6258 2372 6264
rect 3056 6316 3108 6322
rect 3056 6258 3108 6264
rect 2228 6180 2280 6186
rect 2228 6122 2280 6128
rect 1939 6012 2247 6021
rect 1939 6010 1945 6012
rect 2001 6010 2025 6012
rect 2081 6010 2105 6012
rect 2161 6010 2185 6012
rect 2241 6010 2247 6012
rect 2001 5958 2003 6010
rect 2183 5958 2185 6010
rect 1939 5956 1945 5958
rect 2001 5956 2025 5958
rect 2081 5956 2105 5958
rect 2161 5956 2185 5958
rect 2241 5956 2247 5958
rect 1939 5947 2247 5956
rect 2332 5896 2360 6258
rect 2870 6216 2926 6225
rect 2870 6151 2926 6160
rect 2240 5868 2360 5896
rect 2240 5710 2268 5868
rect 2884 5710 2912 6151
rect 3332 6112 3384 6118
rect 3332 6054 3384 6060
rect 1860 5704 1912 5710
rect 1860 5646 1912 5652
rect 2228 5704 2280 5710
rect 2228 5646 2280 5652
rect 2320 5704 2372 5710
rect 2320 5646 2372 5652
rect 2504 5704 2556 5710
rect 2504 5646 2556 5652
rect 2872 5704 2924 5710
rect 2924 5664 3188 5692
rect 2872 5646 2924 5652
rect 1584 5568 1636 5574
rect 1584 5510 1636 5516
rect 1400 5160 1452 5166
rect 1400 5102 1452 5108
rect 1412 3602 1440 5102
rect 1768 5024 1820 5030
rect 1768 4966 1820 4972
rect 1780 4826 1808 4966
rect 1939 4924 2247 4933
rect 1939 4922 1945 4924
rect 2001 4922 2025 4924
rect 2081 4922 2105 4924
rect 2161 4922 2185 4924
rect 2241 4922 2247 4924
rect 2001 4870 2003 4922
rect 2183 4870 2185 4922
rect 1939 4868 1945 4870
rect 2001 4868 2025 4870
rect 2081 4868 2105 4870
rect 2161 4868 2185 4870
rect 2241 4868 2247 4870
rect 1939 4859 2247 4868
rect 1768 4820 1820 4826
rect 1768 4762 1820 4768
rect 2134 4720 2190 4729
rect 2332 4690 2360 5646
rect 2516 5574 2544 5646
rect 2504 5568 2556 5574
rect 2504 5510 2556 5516
rect 2964 5568 3016 5574
rect 2964 5510 3016 5516
rect 2516 5352 2544 5510
rect 2599 5468 2907 5477
rect 2599 5466 2605 5468
rect 2661 5466 2685 5468
rect 2741 5466 2765 5468
rect 2821 5466 2845 5468
rect 2901 5466 2907 5468
rect 2661 5414 2663 5466
rect 2843 5414 2845 5466
rect 2599 5412 2605 5414
rect 2661 5412 2685 5414
rect 2741 5412 2765 5414
rect 2821 5412 2845 5414
rect 2901 5412 2907 5414
rect 2599 5403 2907 5412
rect 2872 5364 2924 5370
rect 2516 5324 2820 5352
rect 2596 5024 2648 5030
rect 2596 4966 2648 4972
rect 2134 4655 2190 4664
rect 2320 4684 2372 4690
rect 1952 4548 2004 4554
rect 1952 4490 2004 4496
rect 1964 4282 1992 4490
rect 2148 4486 2176 4655
rect 2320 4626 2372 4632
rect 2608 4486 2636 4966
rect 2792 4536 2820 5324
rect 2872 5306 2924 5312
rect 2884 4865 2912 5306
rect 2976 5234 3004 5510
rect 3056 5296 3108 5302
rect 3056 5238 3108 5244
rect 2964 5228 3016 5234
rect 2964 5170 3016 5176
rect 2870 4856 2926 4865
rect 3068 4826 3096 5238
rect 3160 4826 3188 5664
rect 3240 5636 3292 5642
rect 3240 5578 3292 5584
rect 3252 5302 3280 5578
rect 3240 5296 3292 5302
rect 3240 5238 3292 5244
rect 2870 4791 2926 4800
rect 3056 4820 3108 4826
rect 3056 4762 3108 4768
rect 3148 4820 3200 4826
rect 3148 4762 3200 4768
rect 3056 4616 3108 4622
rect 3056 4558 3108 4564
rect 2872 4548 2924 4554
rect 2792 4508 2872 4536
rect 2872 4490 2924 4496
rect 2136 4480 2188 4486
rect 2136 4422 2188 4428
rect 2596 4480 2648 4486
rect 2596 4422 2648 4428
rect 1952 4276 2004 4282
rect 1952 4218 2004 4224
rect 1492 4140 1544 4146
rect 1492 4082 1544 4088
rect 1676 4140 1728 4146
rect 2148 4128 2176 4422
rect 2599 4380 2907 4389
rect 2599 4378 2605 4380
rect 2661 4378 2685 4380
rect 2741 4378 2765 4380
rect 2821 4378 2845 4380
rect 2901 4378 2907 4380
rect 2661 4326 2663 4378
rect 2843 4326 2845 4378
rect 2599 4324 2605 4326
rect 2661 4324 2685 4326
rect 2741 4324 2765 4326
rect 2821 4324 2845 4326
rect 2901 4324 2907 4326
rect 2599 4315 2907 4324
rect 2228 4140 2280 4146
rect 2148 4100 2228 4128
rect 1676 4082 1728 4088
rect 2228 4082 2280 4088
rect 2964 4140 3016 4146
rect 2964 4082 3016 4088
rect 1400 3596 1452 3602
rect 1400 3538 1452 3544
rect 1412 3194 1440 3538
rect 1504 3505 1532 4082
rect 1490 3496 1546 3505
rect 1490 3431 1546 3440
rect 1400 3188 1452 3194
rect 1400 3130 1452 3136
rect 20 2848 72 2854
rect 20 2790 72 2796
rect 32 800 60 2790
rect 1688 2774 1716 4082
rect 2320 4072 2372 4078
rect 1766 4040 1822 4049
rect 2320 4014 2372 4020
rect 1766 3975 1768 3984
rect 1820 3975 1822 3984
rect 1768 3946 1820 3952
rect 1860 3936 1912 3942
rect 1860 3878 1912 3884
rect 1872 3194 1900 3878
rect 1939 3836 2247 3845
rect 1939 3834 1945 3836
rect 2001 3834 2025 3836
rect 2081 3834 2105 3836
rect 2161 3834 2185 3836
rect 2241 3834 2247 3836
rect 2001 3782 2003 3834
rect 2183 3782 2185 3834
rect 1939 3780 1945 3782
rect 2001 3780 2025 3782
rect 2081 3780 2105 3782
rect 2161 3780 2185 3782
rect 2241 3780 2247 3782
rect 1939 3771 2247 3780
rect 1860 3188 1912 3194
rect 1860 3130 1912 3136
rect 1768 3052 1820 3058
rect 1768 2994 1820 3000
rect 2044 3052 2096 3058
rect 2044 2994 2096 3000
rect 1596 2746 1716 2774
rect 1596 1902 1624 2746
rect 1780 2650 1808 2994
rect 2056 2961 2084 2994
rect 2042 2952 2098 2961
rect 2042 2887 2098 2896
rect 2332 2854 2360 4014
rect 2872 4004 2924 4010
rect 2872 3946 2924 3952
rect 2412 3936 2464 3942
rect 2412 3878 2464 3884
rect 2504 3936 2556 3942
rect 2504 3878 2556 3884
rect 2424 2938 2452 3878
rect 2516 3738 2544 3878
rect 2884 3738 2912 3946
rect 2504 3732 2556 3738
rect 2504 3674 2556 3680
rect 2872 3732 2924 3738
rect 2872 3674 2924 3680
rect 2976 3602 3004 4082
rect 3068 3602 3096 4558
rect 3252 4486 3280 5238
rect 3344 4486 3372 6054
rect 3436 4622 3464 6820
rect 3516 6724 3568 6730
rect 3516 6666 3568 6672
rect 3528 6322 3556 6666
rect 3620 6390 3648 8871
rect 3712 8294 3740 9522
rect 3884 9512 3936 9518
rect 4160 9512 4212 9518
rect 3936 9472 4160 9500
rect 3884 9454 3936 9460
rect 4160 9454 4212 9460
rect 4344 9512 4396 9518
rect 4344 9454 4396 9460
rect 4436 9512 4488 9518
rect 4436 9454 4488 9460
rect 5816 9512 5868 9518
rect 5816 9454 5868 9460
rect 6368 9512 6420 9518
rect 6368 9454 6420 9460
rect 3917 9276 4225 9285
rect 3917 9274 3923 9276
rect 3979 9274 4003 9276
rect 4059 9274 4083 9276
rect 4139 9274 4163 9276
rect 4219 9274 4225 9276
rect 3979 9222 3981 9274
rect 4161 9222 4163 9274
rect 3917 9220 3923 9222
rect 3979 9220 4003 9222
rect 4059 9220 4083 9222
rect 4139 9220 4163 9222
rect 4219 9220 4225 9222
rect 3917 9211 4225 9220
rect 4068 8968 4120 8974
rect 4068 8910 4120 8916
rect 4080 8498 4108 8910
rect 4356 8906 4384 9454
rect 4344 8900 4396 8906
rect 4344 8842 4396 8848
rect 4252 8832 4304 8838
rect 4252 8774 4304 8780
rect 4068 8492 4120 8498
rect 4068 8434 4120 8440
rect 3700 8288 3752 8294
rect 3700 8230 3752 8236
rect 3712 7954 3740 8230
rect 3917 8188 4225 8197
rect 3917 8186 3923 8188
rect 3979 8186 4003 8188
rect 4059 8186 4083 8188
rect 4139 8186 4163 8188
rect 4219 8186 4225 8188
rect 3979 8134 3981 8186
rect 4161 8134 4163 8186
rect 3917 8132 3923 8134
rect 3979 8132 4003 8134
rect 4059 8132 4083 8134
rect 4139 8132 4163 8134
rect 4219 8132 4225 8134
rect 3917 8123 4225 8132
rect 3884 8016 3936 8022
rect 3884 7958 3936 7964
rect 3700 7948 3752 7954
rect 3700 7890 3752 7896
rect 3700 7744 3752 7750
rect 3700 7686 3752 7692
rect 3792 7744 3844 7750
rect 3792 7686 3844 7692
rect 3608 6384 3660 6390
rect 3608 6326 3660 6332
rect 3516 6316 3568 6322
rect 3516 6258 3568 6264
rect 3528 5710 3556 6258
rect 3608 6112 3660 6118
rect 3608 6054 3660 6060
rect 3516 5704 3568 5710
rect 3516 5646 3568 5652
rect 3528 4758 3556 5646
rect 3516 4752 3568 4758
rect 3516 4694 3568 4700
rect 3424 4616 3476 4622
rect 3424 4558 3476 4564
rect 3240 4480 3292 4486
rect 3240 4422 3292 4428
rect 3332 4480 3384 4486
rect 3332 4422 3384 4428
rect 3240 4004 3292 4010
rect 3240 3946 3292 3952
rect 2964 3596 3016 3602
rect 2964 3538 3016 3544
rect 3056 3596 3108 3602
rect 3056 3538 3108 3544
rect 3068 3398 3096 3538
rect 3252 3534 3280 3946
rect 3436 3738 3464 4558
rect 3620 3738 3648 6054
rect 3712 5778 3740 7686
rect 3804 7410 3832 7686
rect 3792 7404 3844 7410
rect 3792 7346 3844 7352
rect 3896 7188 3924 7958
rect 4264 7342 4292 8774
rect 4448 8294 4476 9454
rect 5172 9444 5224 9450
rect 5172 9386 5224 9392
rect 4577 8732 4885 8741
rect 4577 8730 4583 8732
rect 4639 8730 4663 8732
rect 4719 8730 4743 8732
rect 4799 8730 4823 8732
rect 4879 8730 4885 8732
rect 4639 8678 4641 8730
rect 4821 8678 4823 8730
rect 4577 8676 4583 8678
rect 4639 8676 4663 8678
rect 4719 8676 4743 8678
rect 4799 8676 4823 8678
rect 4879 8676 4885 8678
rect 4577 8667 4885 8676
rect 5080 8560 5132 8566
rect 5080 8502 5132 8508
rect 4436 8288 4488 8294
rect 4436 8230 4488 8236
rect 4988 7948 5040 7954
rect 4988 7890 5040 7896
rect 4436 7880 4488 7886
rect 4356 7840 4436 7868
rect 4356 7546 4384 7840
rect 4436 7822 4488 7828
rect 4436 7744 4488 7750
rect 4436 7686 4488 7692
rect 4344 7540 4396 7546
rect 4344 7482 4396 7488
rect 4344 7404 4396 7410
rect 4344 7346 4396 7352
rect 4252 7336 4304 7342
rect 4252 7278 4304 7284
rect 3804 7160 3924 7188
rect 4252 7200 4304 7206
rect 3700 5772 3752 5778
rect 3700 5714 3752 5720
rect 3700 5228 3752 5234
rect 3700 5170 3752 5176
rect 3712 3890 3740 5170
rect 3804 4146 3832 7160
rect 4252 7142 4304 7148
rect 3917 7100 4225 7109
rect 3917 7098 3923 7100
rect 3979 7098 4003 7100
rect 4059 7098 4083 7100
rect 4139 7098 4163 7100
rect 4219 7098 4225 7100
rect 3979 7046 3981 7098
rect 4161 7046 4163 7098
rect 3917 7044 3923 7046
rect 3979 7044 4003 7046
rect 4059 7044 4083 7046
rect 4139 7044 4163 7046
rect 4219 7044 4225 7046
rect 3917 7035 4225 7044
rect 3884 6928 3936 6934
rect 3884 6870 3936 6876
rect 3896 6322 3924 6870
rect 3976 6792 4028 6798
rect 3976 6734 4028 6740
rect 4068 6792 4120 6798
rect 4068 6734 4120 6740
rect 3988 6322 4016 6734
rect 4080 6662 4108 6734
rect 4068 6656 4120 6662
rect 4068 6598 4120 6604
rect 3884 6316 3936 6322
rect 3884 6258 3936 6264
rect 3976 6316 4028 6322
rect 3976 6258 4028 6264
rect 3896 6225 3924 6258
rect 3882 6216 3938 6225
rect 3882 6151 3938 6160
rect 4080 6118 4108 6598
rect 4068 6112 4120 6118
rect 4068 6054 4120 6060
rect 3917 6012 4225 6021
rect 3917 6010 3923 6012
rect 3979 6010 4003 6012
rect 4059 6010 4083 6012
rect 4139 6010 4163 6012
rect 4219 6010 4225 6012
rect 3979 5958 3981 6010
rect 4161 5958 4163 6010
rect 3917 5956 3923 5958
rect 3979 5956 4003 5958
rect 4059 5956 4083 5958
rect 4139 5956 4163 5958
rect 4219 5956 4225 5958
rect 3917 5947 4225 5956
rect 3882 5808 3938 5817
rect 3882 5743 3938 5752
rect 3896 5166 3924 5743
rect 4264 5710 4292 7142
rect 4356 6118 4384 7346
rect 4344 6112 4396 6118
rect 4344 6054 4396 6060
rect 3976 5704 4028 5710
rect 3976 5646 4028 5652
rect 4068 5704 4120 5710
rect 4160 5704 4212 5710
rect 4068 5646 4120 5652
rect 4158 5672 4160 5681
rect 4252 5704 4304 5710
rect 4212 5672 4214 5681
rect 3884 5160 3936 5166
rect 3884 5102 3936 5108
rect 3988 5030 4016 5646
rect 4080 5370 4108 5646
rect 4252 5646 4304 5652
rect 4158 5607 4214 5616
rect 4160 5568 4212 5574
rect 4160 5510 4212 5516
rect 4068 5364 4120 5370
rect 4068 5306 4120 5312
rect 4172 5098 4200 5510
rect 4264 5302 4292 5646
rect 4252 5296 4304 5302
rect 4252 5238 4304 5244
rect 4252 5160 4304 5166
rect 4252 5102 4304 5108
rect 4160 5092 4212 5098
rect 4160 5034 4212 5040
rect 3976 5024 4028 5030
rect 3976 4966 4028 4972
rect 3917 4924 4225 4933
rect 3917 4922 3923 4924
rect 3979 4922 4003 4924
rect 4059 4922 4083 4924
rect 4139 4922 4163 4924
rect 4219 4922 4225 4924
rect 3979 4870 3981 4922
rect 4161 4870 4163 4922
rect 3917 4868 3923 4870
rect 3979 4868 4003 4870
rect 4059 4868 4083 4870
rect 4139 4868 4163 4870
rect 4219 4868 4225 4870
rect 3917 4859 4225 4868
rect 3976 4820 4028 4826
rect 4264 4808 4292 5102
rect 3976 4762 4028 4768
rect 4172 4780 4292 4808
rect 3988 4214 4016 4762
rect 4068 4616 4120 4622
rect 4066 4584 4068 4593
rect 4120 4584 4122 4593
rect 4066 4519 4122 4528
rect 4068 4480 4120 4486
rect 4068 4422 4120 4428
rect 3976 4208 4028 4214
rect 3976 4150 4028 4156
rect 3792 4140 3844 4146
rect 3792 4082 3844 4088
rect 4080 4010 4108 4422
rect 4172 4282 4200 4780
rect 4252 4480 4304 4486
rect 4252 4422 4304 4428
rect 4160 4276 4212 4282
rect 4160 4218 4212 4224
rect 4068 4004 4120 4010
rect 4068 3946 4120 3952
rect 3712 3862 3832 3890
rect 3424 3732 3476 3738
rect 3424 3674 3476 3680
rect 3608 3732 3660 3738
rect 3608 3674 3660 3680
rect 3700 3732 3752 3738
rect 3700 3674 3752 3680
rect 3332 3664 3384 3670
rect 3332 3606 3384 3612
rect 3240 3528 3292 3534
rect 3240 3470 3292 3476
rect 3056 3392 3108 3398
rect 3056 3334 3108 3340
rect 2599 3292 2907 3301
rect 2599 3290 2605 3292
rect 2661 3290 2685 3292
rect 2741 3290 2765 3292
rect 2821 3290 2845 3292
rect 2901 3290 2907 3292
rect 2661 3238 2663 3290
rect 2843 3238 2845 3290
rect 2599 3236 2605 3238
rect 2661 3236 2685 3238
rect 2741 3236 2765 3238
rect 2821 3236 2845 3238
rect 2901 3236 2907 3238
rect 2599 3227 2907 3236
rect 2780 3120 2832 3126
rect 2780 3062 2832 3068
rect 3238 3088 3294 3097
rect 2424 2910 2636 2938
rect 2608 2854 2636 2910
rect 2320 2848 2372 2854
rect 2320 2790 2372 2796
rect 2596 2848 2648 2854
rect 2596 2790 2648 2796
rect 1939 2748 2247 2757
rect 1939 2746 1945 2748
rect 2001 2746 2025 2748
rect 2081 2746 2105 2748
rect 2161 2746 2185 2748
rect 2241 2746 2247 2748
rect 2001 2694 2003 2746
rect 2183 2694 2185 2746
rect 1939 2692 1945 2694
rect 2001 2692 2025 2694
rect 2081 2692 2105 2694
rect 2161 2692 2185 2694
rect 2241 2692 2247 2694
rect 1939 2683 2247 2692
rect 2792 2650 2820 3062
rect 3238 3023 3294 3032
rect 3252 2922 3280 3023
rect 3240 2916 3292 2922
rect 3240 2858 3292 2864
rect 3344 2774 3372 3606
rect 3712 3584 3740 3674
rect 3620 3556 3740 3584
rect 3424 3460 3476 3466
rect 3424 3402 3476 3408
rect 3252 2746 3372 2774
rect 1768 2644 1820 2650
rect 1768 2586 1820 2592
rect 2504 2644 2556 2650
rect 2504 2586 2556 2592
rect 2780 2644 2832 2650
rect 2780 2586 2832 2592
rect 2516 2553 2544 2586
rect 2502 2544 2558 2553
rect 3252 2514 3280 2746
rect 3436 2666 3464 3402
rect 3620 3058 3648 3556
rect 3804 3398 3832 3862
rect 3917 3836 4225 3845
rect 3917 3834 3923 3836
rect 3979 3834 4003 3836
rect 4059 3834 4083 3836
rect 4139 3834 4163 3836
rect 4219 3834 4225 3836
rect 3979 3782 3981 3834
rect 4161 3782 4163 3834
rect 3917 3780 3923 3782
rect 3979 3780 4003 3782
rect 4059 3780 4083 3782
rect 4139 3780 4163 3782
rect 4219 3780 4225 3782
rect 3917 3771 4225 3780
rect 3974 3632 4030 3641
rect 3896 3590 3974 3618
rect 3896 3534 3924 3590
rect 3974 3567 4030 3576
rect 3884 3528 3936 3534
rect 3884 3470 3936 3476
rect 3988 3454 4200 3482
rect 3988 3398 4016 3454
rect 3792 3392 3844 3398
rect 3792 3334 3844 3340
rect 3884 3392 3936 3398
rect 3884 3334 3936 3340
rect 3976 3392 4028 3398
rect 3976 3334 4028 3340
rect 4068 3392 4120 3398
rect 4068 3334 4120 3340
rect 3896 3074 3924 3334
rect 3608 3052 3660 3058
rect 3608 2994 3660 3000
rect 3712 3046 3924 3074
rect 3344 2638 3464 2666
rect 3620 2650 3648 2994
rect 3608 2644 3660 2650
rect 2502 2479 2558 2488
rect 3240 2508 3292 2514
rect 3240 2450 3292 2456
rect 3344 2446 3372 2638
rect 3608 2586 3660 2592
rect 3332 2440 3384 2446
rect 3424 2440 3476 2446
rect 3332 2382 3384 2388
rect 3422 2408 3424 2417
rect 3476 2408 3478 2417
rect 3056 2372 3108 2378
rect 3422 2343 3478 2352
rect 3056 2314 3108 2320
rect 2599 2204 2907 2213
rect 2599 2202 2605 2204
rect 2661 2202 2685 2204
rect 2741 2202 2765 2204
rect 2821 2202 2845 2204
rect 2901 2202 2907 2204
rect 2661 2150 2663 2202
rect 2843 2150 2845 2202
rect 2599 2148 2605 2150
rect 2661 2148 2685 2150
rect 2741 2148 2765 2150
rect 2821 2148 2845 2150
rect 2901 2148 2907 2150
rect 2599 2139 2907 2148
rect 3068 2038 3096 2314
rect 3516 2304 3568 2310
rect 3516 2246 3568 2252
rect 3056 2032 3108 2038
rect 3056 1974 3108 1980
rect 3528 1970 3556 2246
rect 3516 1964 3568 1970
rect 3516 1906 3568 1912
rect 1584 1896 1636 1902
rect 1584 1838 1636 1844
rect 3712 1766 3740 3046
rect 4080 2938 4108 3334
rect 4172 3194 4200 3454
rect 4160 3188 4212 3194
rect 4160 3130 4212 3136
rect 3804 2910 4108 2938
rect 3804 1902 3832 2910
rect 3917 2748 4225 2757
rect 3917 2746 3923 2748
rect 3979 2746 4003 2748
rect 4059 2746 4083 2748
rect 4139 2746 4163 2748
rect 4219 2746 4225 2748
rect 3979 2694 3981 2746
rect 4161 2694 4163 2746
rect 3917 2692 3923 2694
rect 3979 2692 4003 2694
rect 4059 2692 4083 2694
rect 4139 2692 4163 2694
rect 4219 2692 4225 2694
rect 3917 2683 4225 2692
rect 4264 2378 4292 4422
rect 4356 3126 4384 6054
rect 4448 5234 4476 7686
rect 4577 7644 4885 7653
rect 4577 7642 4583 7644
rect 4639 7642 4663 7644
rect 4719 7642 4743 7644
rect 4799 7642 4823 7644
rect 4879 7642 4885 7644
rect 4639 7590 4641 7642
rect 4821 7590 4823 7642
rect 4577 7588 4583 7590
rect 4639 7588 4663 7590
rect 4719 7588 4743 7590
rect 4799 7588 4823 7590
rect 4879 7588 4885 7590
rect 4577 7579 4885 7588
rect 4620 7404 4672 7410
rect 4620 7346 4672 7352
rect 4896 7404 4948 7410
rect 4896 7346 4948 7352
rect 4528 7336 4580 7342
rect 4528 7278 4580 7284
rect 4540 6934 4568 7278
rect 4528 6928 4580 6934
rect 4528 6870 4580 6876
rect 4540 6798 4568 6870
rect 4632 6798 4660 7346
rect 4908 6866 4936 7346
rect 4896 6860 4948 6866
rect 4896 6802 4948 6808
rect 4528 6792 4580 6798
rect 4528 6734 4580 6740
rect 4620 6792 4672 6798
rect 4620 6734 4672 6740
rect 4577 6556 4885 6565
rect 4577 6554 4583 6556
rect 4639 6554 4663 6556
rect 4719 6554 4743 6556
rect 4799 6554 4823 6556
rect 4879 6554 4885 6556
rect 4639 6502 4641 6554
rect 4821 6502 4823 6554
rect 4577 6500 4583 6502
rect 4639 6500 4663 6502
rect 4719 6500 4743 6502
rect 4799 6500 4823 6502
rect 4879 6500 4885 6502
rect 4577 6491 4885 6500
rect 4712 6452 4764 6458
rect 4712 6394 4764 6400
rect 4526 6352 4582 6361
rect 4526 6287 4528 6296
rect 4580 6287 4582 6296
rect 4528 6258 4580 6264
rect 4620 5908 4672 5914
rect 4620 5850 4672 5856
rect 4632 5556 4660 5850
rect 4724 5710 4752 6394
rect 4804 5772 4856 5778
rect 4856 5732 4936 5760
rect 4804 5714 4856 5720
rect 4712 5704 4764 5710
rect 4712 5646 4764 5652
rect 4804 5568 4856 5574
rect 4632 5528 4804 5556
rect 4804 5510 4856 5516
rect 4908 5522 4936 5732
rect 5000 5710 5028 7890
rect 5092 7886 5120 8502
rect 5080 7880 5132 7886
rect 5078 7848 5080 7857
rect 5132 7848 5134 7857
rect 5078 7783 5134 7792
rect 5080 7744 5132 7750
rect 5080 7686 5132 7692
rect 4988 5704 5040 5710
rect 4988 5646 5040 5652
rect 5092 5522 5120 7686
rect 5184 7206 5212 9386
rect 5828 9178 5856 9454
rect 6276 9376 6328 9382
rect 6276 9318 6328 9324
rect 5895 9276 6203 9285
rect 5895 9274 5901 9276
rect 5957 9274 5981 9276
rect 6037 9274 6061 9276
rect 6117 9274 6141 9276
rect 6197 9274 6203 9276
rect 5957 9222 5959 9274
rect 6139 9222 6141 9274
rect 5895 9220 5901 9222
rect 5957 9220 5981 9222
rect 6037 9220 6061 9222
rect 6117 9220 6141 9222
rect 6197 9220 6203 9222
rect 5895 9211 6203 9220
rect 5816 9172 5868 9178
rect 5816 9114 5868 9120
rect 5724 8900 5776 8906
rect 5724 8842 5776 8848
rect 5264 8832 5316 8838
rect 5264 8774 5316 8780
rect 5276 8616 5304 8774
rect 5356 8628 5408 8634
rect 5276 8588 5356 8616
rect 5356 8570 5408 8576
rect 5264 8288 5316 8294
rect 5264 8230 5316 8236
rect 5276 7478 5304 8230
rect 5368 7954 5396 8570
rect 5632 8492 5684 8498
rect 5632 8434 5684 8440
rect 5540 8424 5592 8430
rect 5540 8366 5592 8372
rect 5448 8288 5500 8294
rect 5448 8230 5500 8236
rect 5356 7948 5408 7954
rect 5356 7890 5408 7896
rect 5264 7472 5316 7478
rect 5264 7414 5316 7420
rect 5264 7336 5316 7342
rect 5264 7278 5316 7284
rect 5172 7200 5224 7206
rect 5172 7142 5224 7148
rect 5172 6656 5224 6662
rect 5172 6598 5224 6604
rect 5184 5953 5212 6598
rect 5170 5944 5226 5953
rect 5170 5879 5226 5888
rect 5184 5710 5212 5879
rect 5172 5704 5224 5710
rect 5172 5646 5224 5652
rect 4908 5494 5120 5522
rect 4577 5468 4885 5477
rect 4577 5466 4583 5468
rect 4639 5466 4663 5468
rect 4719 5466 4743 5468
rect 4799 5466 4823 5468
rect 4879 5466 4885 5468
rect 4639 5414 4641 5466
rect 4821 5414 4823 5466
rect 4577 5412 4583 5414
rect 4639 5412 4663 5414
rect 4719 5412 4743 5414
rect 4799 5412 4823 5414
rect 4879 5412 4885 5414
rect 4577 5403 4885 5412
rect 4986 5400 5042 5409
rect 4620 5364 4672 5370
rect 4620 5306 4672 5312
rect 4712 5364 4764 5370
rect 4712 5306 4764 5312
rect 4908 5358 4986 5386
rect 4436 5228 4488 5234
rect 4436 5170 4488 5176
rect 4448 4690 4476 5170
rect 4632 4865 4660 5306
rect 4618 4856 4674 4865
rect 4618 4791 4674 4800
rect 4436 4684 4488 4690
rect 4436 4626 4488 4632
rect 4528 4616 4580 4622
rect 4632 4604 4660 4791
rect 4580 4576 4660 4604
rect 4528 4558 4580 4564
rect 4724 4486 4752 5306
rect 4804 5228 4856 5234
rect 4804 5170 4856 5176
rect 4816 4729 4844 5170
rect 4802 4720 4858 4729
rect 4802 4655 4858 4664
rect 4908 4554 4936 5358
rect 4986 5335 5042 5344
rect 5092 5098 5120 5494
rect 5170 5128 5226 5137
rect 4988 5092 5040 5098
rect 4988 5034 5040 5040
rect 5080 5092 5132 5098
rect 5170 5063 5226 5072
rect 5080 5034 5132 5040
rect 4896 4548 4948 4554
rect 4896 4490 4948 4496
rect 4528 4480 4580 4486
rect 4448 4440 4528 4468
rect 4448 3534 4476 4440
rect 4528 4422 4580 4428
rect 4712 4480 4764 4486
rect 4712 4422 4764 4428
rect 4577 4380 4885 4389
rect 4577 4378 4583 4380
rect 4639 4378 4663 4380
rect 4719 4378 4743 4380
rect 4799 4378 4823 4380
rect 4879 4378 4885 4380
rect 4639 4326 4641 4378
rect 4821 4326 4823 4378
rect 4577 4324 4583 4326
rect 4639 4324 4663 4326
rect 4719 4324 4743 4326
rect 4799 4324 4823 4326
rect 4879 4324 4885 4326
rect 4577 4315 4885 4324
rect 5000 4146 5028 5034
rect 5078 4992 5134 5001
rect 5078 4927 5134 4936
rect 5092 4690 5120 4927
rect 5184 4826 5212 5063
rect 5276 4865 5304 7278
rect 5368 5574 5396 7890
rect 5460 7342 5488 8230
rect 5552 8022 5580 8366
rect 5540 8016 5592 8022
rect 5540 7958 5592 7964
rect 5644 7868 5672 8434
rect 5736 8090 5764 8842
rect 5828 8634 5856 9114
rect 5816 8628 5868 8634
rect 5816 8570 5868 8576
rect 5816 8356 5868 8362
rect 5816 8298 5868 8304
rect 5724 8084 5776 8090
rect 5828 8072 5856 8298
rect 5895 8188 6203 8197
rect 5895 8186 5901 8188
rect 5957 8186 5981 8188
rect 6037 8186 6061 8188
rect 6117 8186 6141 8188
rect 6197 8186 6203 8188
rect 5957 8134 5959 8186
rect 6139 8134 6141 8186
rect 5895 8132 5901 8134
rect 5957 8132 5981 8134
rect 6037 8132 6061 8134
rect 6117 8132 6141 8134
rect 6197 8132 6203 8134
rect 5895 8123 6203 8132
rect 5828 8044 6040 8072
rect 5724 8026 5776 8032
rect 5906 7984 5962 7993
rect 5906 7919 5962 7928
rect 5552 7840 5672 7868
rect 5552 7342 5580 7840
rect 5920 7410 5948 7919
rect 6012 7818 6040 8044
rect 6184 8016 6236 8022
rect 6184 7958 6236 7964
rect 6196 7818 6224 7958
rect 6000 7812 6052 7818
rect 6000 7754 6052 7760
rect 6092 7812 6144 7818
rect 6092 7754 6144 7760
rect 6184 7812 6236 7818
rect 6184 7754 6236 7760
rect 5908 7404 5960 7410
rect 5736 7364 5908 7392
rect 5448 7336 5500 7342
rect 5448 7278 5500 7284
rect 5540 7336 5592 7342
rect 5540 7278 5592 7284
rect 5630 7304 5686 7313
rect 5460 6662 5488 7278
rect 5630 7239 5686 7248
rect 5540 6928 5592 6934
rect 5540 6870 5592 6876
rect 5448 6656 5500 6662
rect 5448 6598 5500 6604
rect 5552 5914 5580 6870
rect 5644 6390 5672 7239
rect 5736 6934 5764 7364
rect 5908 7346 5960 7352
rect 6104 7313 6132 7754
rect 6090 7304 6146 7313
rect 6288 7290 6316 9318
rect 6380 8401 6408 9454
rect 6366 8392 6422 8401
rect 6366 8327 6422 8336
rect 6368 8288 6420 8294
rect 6368 8230 6420 8236
rect 6380 8090 6408 8230
rect 6368 8084 6420 8090
rect 6368 8026 6420 8032
rect 6366 7848 6422 7857
rect 6366 7783 6422 7792
rect 6380 7750 6408 7783
rect 6368 7744 6420 7750
rect 6368 7686 6420 7692
rect 6380 7410 6408 7686
rect 6472 7426 6500 9522
rect 6920 9512 6972 9518
rect 6920 9454 6972 9460
rect 6555 8732 6863 8741
rect 6555 8730 6561 8732
rect 6617 8730 6641 8732
rect 6697 8730 6721 8732
rect 6777 8730 6801 8732
rect 6857 8730 6863 8732
rect 6617 8678 6619 8730
rect 6799 8678 6801 8730
rect 6555 8676 6561 8678
rect 6617 8676 6641 8678
rect 6697 8676 6721 8678
rect 6777 8676 6801 8678
rect 6857 8676 6863 8678
rect 6555 8667 6863 8676
rect 6736 8560 6788 8566
rect 6736 8502 6788 8508
rect 6644 8492 6696 8498
rect 6644 8434 6696 8440
rect 6552 8356 6604 8362
rect 6552 8298 6604 8304
rect 6564 7954 6592 8298
rect 6552 7948 6604 7954
rect 6552 7890 6604 7896
rect 6656 7886 6684 8434
rect 6748 8090 6776 8502
rect 6736 8084 6788 8090
rect 6736 8026 6788 8032
rect 6644 7880 6696 7886
rect 6644 7822 6696 7828
rect 6555 7644 6863 7653
rect 6555 7642 6561 7644
rect 6617 7642 6641 7644
rect 6697 7642 6721 7644
rect 6777 7642 6801 7644
rect 6857 7642 6863 7644
rect 6617 7590 6619 7642
rect 6799 7590 6801 7642
rect 6555 7588 6561 7590
rect 6617 7588 6641 7590
rect 6697 7588 6721 7590
rect 6777 7588 6801 7590
rect 6857 7588 6863 7590
rect 6555 7579 6863 7588
rect 6472 7410 6868 7426
rect 6368 7404 6420 7410
rect 6368 7346 6420 7352
rect 6472 7404 6880 7410
rect 6472 7398 6828 7404
rect 6288 7262 6408 7290
rect 6090 7239 6146 7248
rect 6276 7200 6328 7206
rect 6276 7142 6328 7148
rect 5895 7100 6203 7109
rect 5895 7098 5901 7100
rect 5957 7098 5981 7100
rect 6037 7098 6061 7100
rect 6117 7098 6141 7100
rect 6197 7098 6203 7100
rect 5957 7046 5959 7098
rect 6139 7046 6141 7098
rect 5895 7044 5901 7046
rect 5957 7044 5981 7046
rect 6037 7044 6061 7046
rect 6117 7044 6141 7046
rect 6197 7044 6203 7046
rect 5895 7035 6203 7044
rect 5724 6928 5776 6934
rect 5724 6870 5776 6876
rect 5816 6928 5868 6934
rect 5816 6870 5868 6876
rect 5724 6792 5776 6798
rect 5724 6734 5776 6740
rect 5632 6384 5684 6390
rect 5632 6326 5684 6332
rect 5736 6322 5764 6734
rect 5828 6390 5856 6870
rect 6184 6792 6236 6798
rect 6184 6734 6236 6740
rect 6196 6390 6224 6734
rect 5816 6384 5868 6390
rect 5816 6326 5868 6332
rect 6184 6384 6236 6390
rect 6184 6326 6236 6332
rect 5724 6316 5776 6322
rect 5724 6258 5776 6264
rect 5540 5908 5592 5914
rect 5540 5850 5592 5856
rect 5828 5846 5856 6326
rect 5895 6012 6203 6021
rect 5895 6010 5901 6012
rect 5957 6010 5981 6012
rect 6037 6010 6061 6012
rect 6117 6010 6141 6012
rect 6197 6010 6203 6012
rect 5957 5958 5959 6010
rect 6139 5958 6141 6010
rect 5895 5956 5901 5958
rect 5957 5956 5981 5958
rect 6037 5956 6061 5958
rect 6117 5956 6141 5958
rect 6197 5956 6203 5958
rect 5895 5947 6203 5956
rect 6000 5908 6052 5914
rect 6000 5850 6052 5856
rect 5816 5840 5868 5846
rect 5868 5800 5948 5828
rect 5816 5782 5868 5788
rect 5448 5772 5500 5778
rect 5632 5772 5684 5778
rect 5448 5714 5500 5720
rect 5552 5732 5632 5760
rect 5356 5568 5408 5574
rect 5356 5510 5408 5516
rect 5356 5364 5408 5370
rect 5356 5306 5408 5312
rect 5368 5234 5396 5306
rect 5460 5302 5488 5714
rect 5552 5681 5580 5732
rect 5632 5714 5684 5720
rect 5538 5672 5594 5681
rect 5538 5607 5594 5616
rect 5448 5296 5500 5302
rect 5448 5238 5500 5244
rect 5356 5228 5408 5234
rect 5356 5170 5408 5176
rect 5356 5024 5408 5030
rect 5356 4966 5408 4972
rect 5448 5024 5500 5030
rect 5448 4966 5500 4972
rect 5262 4856 5318 4865
rect 5172 4820 5224 4826
rect 5262 4791 5318 4800
rect 5172 4762 5224 4768
rect 5080 4684 5132 4690
rect 5080 4626 5132 4632
rect 5276 4457 5304 4791
rect 5262 4448 5318 4457
rect 5262 4383 5318 4392
rect 4988 4140 5040 4146
rect 4988 4082 5040 4088
rect 4528 4072 4580 4078
rect 4528 4014 4580 4020
rect 4540 3534 4568 4014
rect 4620 3732 4672 3738
rect 4620 3674 4672 3680
rect 4632 3534 4660 3674
rect 5000 3534 5028 4082
rect 5172 3664 5224 3670
rect 5170 3632 5172 3641
rect 5224 3632 5226 3641
rect 5170 3567 5226 3576
rect 4436 3528 4488 3534
rect 4436 3470 4488 3476
rect 4528 3528 4580 3534
rect 4528 3470 4580 3476
rect 4620 3528 4672 3534
rect 4620 3470 4672 3476
rect 4988 3528 5040 3534
rect 5172 3528 5224 3534
rect 5040 3476 5120 3482
rect 4988 3470 5120 3476
rect 5172 3470 5224 3476
rect 5264 3528 5316 3534
rect 5264 3470 5316 3476
rect 4632 3398 4660 3470
rect 5000 3454 5120 3470
rect 4620 3392 4672 3398
rect 4620 3334 4672 3340
rect 4988 3392 5040 3398
rect 4988 3334 5040 3340
rect 4577 3292 4885 3301
rect 4577 3290 4583 3292
rect 4639 3290 4663 3292
rect 4719 3290 4743 3292
rect 4799 3290 4823 3292
rect 4879 3290 4885 3292
rect 4639 3238 4641 3290
rect 4821 3238 4823 3290
rect 4577 3236 4583 3238
rect 4639 3236 4663 3238
rect 4719 3236 4743 3238
rect 4799 3236 4823 3238
rect 4879 3236 4885 3238
rect 4577 3227 4885 3236
rect 5000 3194 5028 3334
rect 4896 3188 4948 3194
rect 4896 3130 4948 3136
rect 4988 3188 5040 3194
rect 4988 3130 5040 3136
rect 4344 3120 4396 3126
rect 4344 3062 4396 3068
rect 4908 3074 4936 3130
rect 5092 3074 5120 3454
rect 4908 3046 5120 3074
rect 4988 2984 5040 2990
rect 5184 2938 5212 3470
rect 4988 2926 5040 2932
rect 5000 2650 5028 2926
rect 5092 2910 5212 2938
rect 4988 2644 5040 2650
rect 4988 2586 5040 2592
rect 5092 2553 5120 2910
rect 5172 2848 5224 2854
rect 5172 2790 5224 2796
rect 5078 2544 5134 2553
rect 5078 2479 5134 2488
rect 5184 2378 5212 2790
rect 5276 2446 5304 3470
rect 5264 2440 5316 2446
rect 5264 2382 5316 2388
rect 4252 2372 4304 2378
rect 4252 2314 4304 2320
rect 5172 2372 5224 2378
rect 5172 2314 5224 2320
rect 4577 2204 4885 2213
rect 4577 2202 4583 2204
rect 4639 2202 4663 2204
rect 4719 2202 4743 2204
rect 4799 2202 4823 2204
rect 4879 2202 4885 2204
rect 4639 2150 4641 2202
rect 4821 2150 4823 2202
rect 4577 2148 4583 2150
rect 4639 2148 4663 2150
rect 4719 2148 4743 2150
rect 4799 2148 4823 2150
rect 4879 2148 4885 2150
rect 4577 2139 4885 2148
rect 5368 2038 5396 4966
rect 5460 4758 5488 4966
rect 5448 4752 5500 4758
rect 5448 4694 5500 4700
rect 5448 4548 5500 4554
rect 5448 4490 5500 4496
rect 5460 3108 5488 4490
rect 5552 4486 5580 5607
rect 5632 5568 5684 5574
rect 5632 5510 5684 5516
rect 5644 5234 5672 5510
rect 5724 5296 5776 5302
rect 5724 5238 5776 5244
rect 5632 5228 5684 5234
rect 5632 5170 5684 5176
rect 5644 5001 5672 5170
rect 5630 4992 5686 5001
rect 5630 4927 5686 4936
rect 5632 4616 5684 4622
rect 5632 4558 5684 4564
rect 5540 4480 5592 4486
rect 5540 4422 5592 4428
rect 5552 4214 5580 4422
rect 5540 4208 5592 4214
rect 5540 4150 5592 4156
rect 5644 4146 5672 4558
rect 5632 4140 5684 4146
rect 5632 4082 5684 4088
rect 5540 3936 5592 3942
rect 5540 3878 5592 3884
rect 5632 3936 5684 3942
rect 5632 3878 5684 3884
rect 5552 3738 5580 3878
rect 5540 3732 5592 3738
rect 5540 3674 5592 3680
rect 5644 3194 5672 3878
rect 5632 3188 5684 3194
rect 5632 3130 5684 3136
rect 5540 3120 5592 3126
rect 5460 3080 5540 3108
rect 5540 3062 5592 3068
rect 5552 2446 5580 3062
rect 5632 2984 5684 2990
rect 5632 2926 5684 2932
rect 5644 2650 5672 2926
rect 5632 2644 5684 2650
rect 5632 2586 5684 2592
rect 5540 2440 5592 2446
rect 5632 2440 5684 2446
rect 5540 2382 5592 2388
rect 5630 2408 5632 2417
rect 5684 2408 5686 2417
rect 5630 2343 5686 2352
rect 5736 2038 5764 5238
rect 5816 5092 5868 5098
rect 5816 5034 5868 5040
rect 5828 4672 5856 5034
rect 5920 5012 5948 5800
rect 6012 5114 6040 5850
rect 6288 5658 6316 7142
rect 6380 7002 6408 7262
rect 6368 6996 6420 7002
rect 6368 6938 6420 6944
rect 6472 6934 6500 7398
rect 6828 7346 6880 7352
rect 6736 7336 6788 7342
rect 6736 7278 6788 7284
rect 6748 7002 6776 7278
rect 6736 6996 6788 7002
rect 6736 6938 6788 6944
rect 6460 6928 6512 6934
rect 6460 6870 6512 6876
rect 6932 6798 6960 9454
rect 7104 9376 7156 9382
rect 7104 9318 7156 9324
rect 7012 7744 7064 7750
rect 7012 7686 7064 7692
rect 7024 6798 7052 7686
rect 7116 7478 7144 9318
rect 7392 8974 7420 9522
rect 7380 8968 7432 8974
rect 7380 8910 7432 8916
rect 7288 8424 7340 8430
rect 7392 8412 7420 8910
rect 7576 8650 7604 9522
rect 8392 9376 8444 9382
rect 8392 9318 8444 9324
rect 7873 9276 8181 9285
rect 7873 9274 7879 9276
rect 7935 9274 7959 9276
rect 8015 9274 8039 9276
rect 8095 9274 8119 9276
rect 8175 9274 8181 9276
rect 7935 9222 7937 9274
rect 8117 9222 8119 9274
rect 7873 9220 7879 9222
rect 7935 9220 7959 9222
rect 8015 9220 8039 9222
rect 8095 9220 8119 9222
rect 8175 9220 8181 9222
rect 7873 9211 8181 9220
rect 7656 8968 7708 8974
rect 7656 8910 7708 8916
rect 8300 8968 8352 8974
rect 8404 8922 8432 9318
rect 8352 8916 8432 8922
rect 8300 8910 8432 8916
rect 7340 8384 7420 8412
rect 7484 8622 7604 8650
rect 7668 8634 7696 8910
rect 8312 8894 8432 8910
rect 7748 8832 7800 8838
rect 7748 8774 7800 8780
rect 7656 8628 7708 8634
rect 7288 8366 7340 8372
rect 7196 8288 7248 8294
rect 7196 8230 7248 8236
rect 7208 8090 7236 8230
rect 7196 8084 7248 8090
rect 7196 8026 7248 8032
rect 7196 7540 7248 7546
rect 7196 7482 7248 7488
rect 7104 7472 7156 7478
rect 7104 7414 7156 7420
rect 6460 6792 6512 6798
rect 6460 6734 6512 6740
rect 6920 6792 6972 6798
rect 6920 6734 6972 6740
rect 7012 6792 7064 6798
rect 7064 6752 7144 6780
rect 7012 6734 7064 6740
rect 6472 6662 6500 6734
rect 6460 6656 6512 6662
rect 6460 6598 6512 6604
rect 6555 6556 6863 6565
rect 6555 6554 6561 6556
rect 6617 6554 6641 6556
rect 6697 6554 6721 6556
rect 6777 6554 6801 6556
rect 6857 6554 6863 6556
rect 6617 6502 6619 6554
rect 6799 6502 6801 6554
rect 6555 6500 6561 6502
rect 6617 6500 6641 6502
rect 6697 6500 6721 6502
rect 6777 6500 6801 6502
rect 6857 6500 6863 6502
rect 6555 6491 6863 6500
rect 6932 6322 6960 6734
rect 7012 6656 7064 6662
rect 7012 6598 7064 6604
rect 6368 6316 6420 6322
rect 6368 6258 6420 6264
rect 6920 6316 6972 6322
rect 6920 6258 6972 6264
rect 6196 5630 6316 5658
rect 6196 5234 6224 5630
rect 6276 5568 6328 5574
rect 6276 5510 6328 5516
rect 6184 5228 6236 5234
rect 6184 5170 6236 5176
rect 6090 5128 6146 5137
rect 6012 5086 6090 5114
rect 6090 5063 6146 5072
rect 6000 5024 6052 5030
rect 5920 4984 6000 5012
rect 6000 4966 6052 4972
rect 5895 4924 6203 4933
rect 5895 4922 5901 4924
rect 5957 4922 5981 4924
rect 6037 4922 6061 4924
rect 6117 4922 6141 4924
rect 6197 4922 6203 4924
rect 5957 4870 5959 4922
rect 6139 4870 6141 4922
rect 5895 4868 5901 4870
rect 5957 4868 5981 4870
rect 6037 4868 6061 4870
rect 6117 4868 6141 4870
rect 6197 4868 6203 4870
rect 5895 4859 6203 4868
rect 6184 4684 6236 4690
rect 5828 4644 6184 4672
rect 6184 4626 6236 4632
rect 5998 4584 6054 4593
rect 6288 4570 6316 5510
rect 6380 5370 6408 6258
rect 6460 6112 6512 6118
rect 6460 6054 6512 6060
rect 6472 5846 6500 6054
rect 7024 5914 7052 6598
rect 7012 5908 7064 5914
rect 7012 5850 7064 5856
rect 6460 5840 6512 5846
rect 6460 5782 6512 5788
rect 6460 5704 6512 5710
rect 6460 5646 6512 5652
rect 6920 5704 6972 5710
rect 6920 5646 6972 5652
rect 7012 5704 7064 5710
rect 7012 5646 7064 5652
rect 6368 5364 6420 5370
rect 6368 5306 6420 5312
rect 6054 4542 6316 4570
rect 5998 4519 6054 4528
rect 6012 4486 6040 4519
rect 5908 4480 5960 4486
rect 5908 4422 5960 4428
rect 6000 4480 6052 4486
rect 6000 4422 6052 4428
rect 6184 4480 6236 4486
rect 6184 4422 6236 4428
rect 5920 4282 5948 4422
rect 5908 4276 5960 4282
rect 5908 4218 5960 4224
rect 6196 4078 6224 4422
rect 6276 4140 6328 4146
rect 6276 4082 6328 4088
rect 6184 4072 6236 4078
rect 6184 4014 6236 4020
rect 5895 3836 6203 3845
rect 5895 3834 5901 3836
rect 5957 3834 5981 3836
rect 6037 3834 6061 3836
rect 6117 3834 6141 3836
rect 6197 3834 6203 3836
rect 5957 3782 5959 3834
rect 6139 3782 6141 3834
rect 5895 3780 5901 3782
rect 5957 3780 5981 3782
rect 6037 3780 6061 3782
rect 6117 3780 6141 3782
rect 6197 3780 6203 3782
rect 5895 3771 6203 3780
rect 6288 3720 6316 4082
rect 6380 3942 6408 5306
rect 6472 5273 6500 5646
rect 6555 5468 6863 5477
rect 6555 5466 6561 5468
rect 6617 5466 6641 5468
rect 6697 5466 6721 5468
rect 6777 5466 6801 5468
rect 6857 5466 6863 5468
rect 6617 5414 6619 5466
rect 6799 5414 6801 5466
rect 6555 5412 6561 5414
rect 6617 5412 6641 5414
rect 6697 5412 6721 5414
rect 6777 5412 6801 5414
rect 6857 5412 6863 5414
rect 6555 5403 6863 5412
rect 6932 5370 6960 5646
rect 6920 5364 6972 5370
rect 6920 5306 6972 5312
rect 6458 5264 6514 5273
rect 6458 5199 6514 5208
rect 6644 5228 6696 5234
rect 6472 4826 6500 5199
rect 6644 5170 6696 5176
rect 6656 5137 6684 5170
rect 6642 5128 6698 5137
rect 6642 5063 6644 5072
rect 6696 5063 6698 5072
rect 6644 5034 6696 5040
rect 6736 5024 6788 5030
rect 6736 4966 6788 4972
rect 6748 4826 6776 4966
rect 7024 4826 7052 5646
rect 7116 5556 7144 6752
rect 7208 5710 7236 7482
rect 7300 6322 7328 8366
rect 7380 8016 7432 8022
rect 7380 7958 7432 7964
rect 7392 6798 7420 7958
rect 7484 7818 7512 8622
rect 7656 8570 7708 8576
rect 7564 8492 7616 8498
rect 7564 8434 7616 8440
rect 7576 8090 7604 8434
rect 7564 8084 7616 8090
rect 7564 8026 7616 8032
rect 7760 8022 7788 8774
rect 8404 8294 8432 8894
rect 8533 8732 8841 8741
rect 8533 8730 8539 8732
rect 8595 8730 8619 8732
rect 8675 8730 8699 8732
rect 8755 8730 8779 8732
rect 8835 8730 8841 8732
rect 8595 8678 8597 8730
rect 8777 8678 8779 8730
rect 8533 8676 8539 8678
rect 8595 8676 8619 8678
rect 8675 8676 8699 8678
rect 8755 8676 8779 8678
rect 8835 8676 8841 8678
rect 8533 8667 8841 8676
rect 8392 8288 8444 8294
rect 8392 8230 8444 8236
rect 8668 8288 8720 8294
rect 8668 8230 8720 8236
rect 7873 8188 8181 8197
rect 7873 8186 7879 8188
rect 7935 8186 7959 8188
rect 8015 8186 8039 8188
rect 8095 8186 8119 8188
rect 8175 8186 8181 8188
rect 7935 8134 7937 8186
rect 8117 8134 8119 8186
rect 7873 8132 7879 8134
rect 7935 8132 7959 8134
rect 8015 8132 8039 8134
rect 8095 8132 8119 8134
rect 8175 8132 8181 8134
rect 7873 8123 8181 8132
rect 7656 8016 7708 8022
rect 7562 7984 7618 7993
rect 7656 7958 7708 7964
rect 7748 8016 7800 8022
rect 7748 7958 7800 7964
rect 8114 7984 8170 7993
rect 7562 7919 7564 7928
rect 7616 7919 7618 7928
rect 7564 7890 7616 7896
rect 7668 7834 7696 7958
rect 8114 7919 8170 7928
rect 8024 7880 8076 7886
rect 7668 7828 8024 7834
rect 7668 7822 8076 7828
rect 7472 7812 7524 7818
rect 7472 7754 7524 7760
rect 7564 7812 7616 7818
rect 7668 7806 8064 7822
rect 7564 7754 7616 7760
rect 7472 7472 7524 7478
rect 7472 7414 7524 7420
rect 7484 6866 7512 7414
rect 7472 6860 7524 6866
rect 7472 6802 7524 6808
rect 7380 6792 7432 6798
rect 7380 6734 7432 6740
rect 7392 6458 7420 6734
rect 7472 6656 7524 6662
rect 7472 6598 7524 6604
rect 7484 6458 7512 6598
rect 7380 6452 7432 6458
rect 7380 6394 7432 6400
rect 7472 6452 7524 6458
rect 7472 6394 7524 6400
rect 7288 6316 7340 6322
rect 7288 6258 7340 6264
rect 7288 6112 7340 6118
rect 7288 6054 7340 6060
rect 7196 5704 7248 5710
rect 7196 5646 7248 5652
rect 7116 5528 7236 5556
rect 6460 4820 6512 4826
rect 6460 4762 6512 4768
rect 6736 4820 6788 4826
rect 6736 4762 6788 4768
rect 7012 4820 7064 4826
rect 7012 4762 7064 4768
rect 6458 4720 6514 4729
rect 6458 4655 6514 4664
rect 6472 4622 6500 4655
rect 7208 4622 7236 5528
rect 6460 4616 6512 4622
rect 6460 4558 6512 4564
rect 7012 4616 7064 4622
rect 7012 4558 7064 4564
rect 7196 4616 7248 4622
rect 7196 4558 7248 4564
rect 6828 4480 6880 4486
rect 6880 4440 6960 4468
rect 6828 4422 6880 4428
rect 6555 4380 6863 4389
rect 6555 4378 6561 4380
rect 6617 4378 6641 4380
rect 6697 4378 6721 4380
rect 6777 4378 6801 4380
rect 6857 4378 6863 4380
rect 6617 4326 6619 4378
rect 6799 4326 6801 4378
rect 6555 4324 6561 4326
rect 6617 4324 6641 4326
rect 6697 4324 6721 4326
rect 6777 4324 6801 4326
rect 6857 4324 6863 4326
rect 6555 4315 6863 4324
rect 6932 4162 6960 4440
rect 7024 4321 7052 4558
rect 7104 4548 7156 4554
rect 7104 4490 7156 4496
rect 7010 4312 7066 4321
rect 7116 4282 7144 4490
rect 7010 4247 7066 4256
rect 7104 4276 7156 4282
rect 7104 4218 7156 4224
rect 6932 4146 7144 4162
rect 6828 4140 6880 4146
rect 6932 4140 7156 4146
rect 6932 4134 7104 4140
rect 6828 4082 6880 4088
rect 7104 4082 7156 4088
rect 6736 4004 6788 4010
rect 6736 3946 6788 3952
rect 6368 3936 6420 3942
rect 6368 3878 6420 3884
rect 6288 3692 6500 3720
rect 6276 3460 6328 3466
rect 6276 3402 6328 3408
rect 5908 3052 5960 3058
rect 5908 2994 5960 3000
rect 5816 2916 5868 2922
rect 5920 2904 5948 2994
rect 5868 2876 5948 2904
rect 5816 2858 5868 2864
rect 5828 2446 5856 2858
rect 5895 2748 6203 2757
rect 5895 2746 5901 2748
rect 5957 2746 5981 2748
rect 6037 2746 6061 2748
rect 6117 2746 6141 2748
rect 6197 2746 6203 2748
rect 5957 2694 5959 2746
rect 6139 2694 6141 2746
rect 5895 2692 5901 2694
rect 5957 2692 5981 2694
rect 6037 2692 6061 2694
rect 6117 2692 6141 2694
rect 6197 2692 6203 2694
rect 5895 2683 6203 2692
rect 6288 2650 6316 3402
rect 6368 2848 6420 2854
rect 6368 2790 6420 2796
rect 5908 2644 5960 2650
rect 5908 2586 5960 2592
rect 6276 2644 6328 2650
rect 6276 2586 6328 2592
rect 5920 2446 5948 2586
rect 6380 2514 6408 2790
rect 6472 2582 6500 3692
rect 6748 3602 6776 3946
rect 6736 3596 6788 3602
rect 6736 3538 6788 3544
rect 6840 3482 6868 4082
rect 7012 4004 7064 4010
rect 7012 3946 7064 3952
rect 7024 3516 7052 3946
rect 7208 3942 7236 4558
rect 7196 3936 7248 3942
rect 7196 3878 7248 3884
rect 7104 3528 7156 3534
rect 7024 3488 7104 3516
rect 6840 3454 6960 3482
rect 7104 3470 7156 3476
rect 7300 3466 7328 6054
rect 7576 5914 7604 7754
rect 8128 7750 8156 7919
rect 8404 7886 8432 8230
rect 8392 7880 8444 7886
rect 8392 7822 8444 7828
rect 8300 7812 8352 7818
rect 8300 7754 8352 7760
rect 8116 7744 8168 7750
rect 8168 7704 8248 7732
rect 8116 7686 8168 7692
rect 7840 7540 7892 7546
rect 7840 7482 7892 7488
rect 7852 7274 7880 7482
rect 8220 7478 8248 7704
rect 8312 7546 8340 7754
rect 8300 7540 8352 7546
rect 8300 7482 8352 7488
rect 8208 7472 8260 7478
rect 8208 7414 8260 7420
rect 7840 7268 7892 7274
rect 7840 7210 7892 7216
rect 7748 7200 7800 7206
rect 7748 7142 7800 7148
rect 7760 6746 7788 7142
rect 7873 7100 8181 7109
rect 7873 7098 7879 7100
rect 7935 7098 7959 7100
rect 8015 7098 8039 7100
rect 8095 7098 8119 7100
rect 8175 7098 8181 7100
rect 7935 7046 7937 7098
rect 8117 7046 8119 7098
rect 7873 7044 7879 7046
rect 7935 7044 7959 7046
rect 8015 7044 8039 7046
rect 8095 7044 8119 7046
rect 8175 7044 8181 7046
rect 7873 7035 8181 7044
rect 8220 6984 8248 7414
rect 8300 7404 8352 7410
rect 8300 7346 8352 7352
rect 8128 6956 8248 6984
rect 7760 6718 7880 6746
rect 8128 6730 8156 6956
rect 8312 6866 8340 7346
rect 8404 7274 8432 7822
rect 8680 7750 8708 8230
rect 8668 7744 8720 7750
rect 8668 7686 8720 7692
rect 8533 7644 8841 7653
rect 8533 7642 8539 7644
rect 8595 7642 8619 7644
rect 8675 7642 8699 7644
rect 8755 7642 8779 7644
rect 8835 7642 8841 7644
rect 8595 7590 8597 7642
rect 8777 7590 8779 7642
rect 8533 7588 8539 7590
rect 8595 7588 8619 7590
rect 8675 7588 8699 7590
rect 8755 7588 8779 7590
rect 8835 7588 8841 7590
rect 8533 7579 8841 7588
rect 9034 7576 9090 7585
rect 9034 7511 9090 7520
rect 8392 7268 8444 7274
rect 8392 7210 8444 7216
rect 8404 7002 8432 7210
rect 8484 7200 8536 7206
rect 8484 7142 8536 7148
rect 8392 6996 8444 7002
rect 8392 6938 8444 6944
rect 8300 6860 8352 6866
rect 8300 6802 8352 6808
rect 8208 6792 8260 6798
rect 8404 6746 8432 6938
rect 8208 6734 8260 6740
rect 7656 6656 7708 6662
rect 7656 6598 7708 6604
rect 7748 6656 7800 6662
rect 7748 6598 7800 6604
rect 7564 5908 7616 5914
rect 7564 5850 7616 5856
rect 7668 5794 7696 6598
rect 7760 5914 7788 6598
rect 7852 6100 7880 6718
rect 8116 6724 8168 6730
rect 8116 6666 8168 6672
rect 7932 6112 7984 6118
rect 7852 6072 7932 6100
rect 7932 6054 7984 6060
rect 7873 6012 8181 6021
rect 7873 6010 7879 6012
rect 7935 6010 7959 6012
rect 8015 6010 8039 6012
rect 8095 6010 8119 6012
rect 8175 6010 8181 6012
rect 7935 5958 7937 6010
rect 8117 5958 8119 6010
rect 7873 5956 7879 5958
rect 7935 5956 7959 5958
rect 8015 5956 8039 5958
rect 8095 5956 8119 5958
rect 8175 5956 8181 5958
rect 7873 5947 8181 5956
rect 8220 5914 8248 6734
rect 8312 6718 8432 6746
rect 7748 5908 7800 5914
rect 7748 5850 7800 5856
rect 8208 5908 8260 5914
rect 8208 5850 8260 5856
rect 7576 5766 7696 5794
rect 7472 5568 7524 5574
rect 7472 5510 7524 5516
rect 7484 5370 7512 5510
rect 7472 5364 7524 5370
rect 7472 5306 7524 5312
rect 7484 4826 7512 5306
rect 7576 5302 7604 5766
rect 7656 5704 7708 5710
rect 7656 5646 7708 5652
rect 8208 5704 8260 5710
rect 8208 5646 8260 5652
rect 7564 5296 7616 5302
rect 7564 5238 7616 5244
rect 7668 5166 7696 5646
rect 8220 5234 8248 5646
rect 8312 5302 8340 6718
rect 8392 6656 8444 6662
rect 8496 6644 8524 7142
rect 8944 6860 8996 6866
rect 8944 6802 8996 6808
rect 8444 6616 8524 6644
rect 8392 6598 8444 6604
rect 8404 5846 8432 6598
rect 8533 6556 8841 6565
rect 8533 6554 8539 6556
rect 8595 6554 8619 6556
rect 8675 6554 8699 6556
rect 8755 6554 8779 6556
rect 8835 6554 8841 6556
rect 8595 6502 8597 6554
rect 8777 6502 8779 6554
rect 8533 6500 8539 6502
rect 8595 6500 8619 6502
rect 8675 6500 8699 6502
rect 8755 6500 8779 6502
rect 8835 6500 8841 6502
rect 8533 6491 8841 6500
rect 8956 6118 8984 6802
rect 9048 6798 9076 7511
rect 9036 6792 9088 6798
rect 9036 6734 9088 6740
rect 8944 6112 8996 6118
rect 8944 6054 8996 6060
rect 8392 5840 8444 5846
rect 8392 5782 8444 5788
rect 8392 5704 8444 5710
rect 8392 5646 8444 5652
rect 8300 5296 8352 5302
rect 8300 5238 8352 5244
rect 8404 5234 8432 5646
rect 8533 5468 8841 5477
rect 8533 5466 8539 5468
rect 8595 5466 8619 5468
rect 8675 5466 8699 5468
rect 8755 5466 8779 5468
rect 8835 5466 8841 5468
rect 8595 5414 8597 5466
rect 8777 5414 8779 5466
rect 8533 5412 8539 5414
rect 8595 5412 8619 5414
rect 8675 5412 8699 5414
rect 8755 5412 8779 5414
rect 8835 5412 8841 5414
rect 8533 5403 8841 5412
rect 8208 5228 8260 5234
rect 8208 5170 8260 5176
rect 8392 5228 8444 5234
rect 8392 5170 8444 5176
rect 7656 5160 7708 5166
rect 7656 5102 7708 5108
rect 7748 5160 7800 5166
rect 7748 5102 7800 5108
rect 7564 5024 7616 5030
rect 7564 4966 7616 4972
rect 7472 4820 7524 4826
rect 7472 4762 7524 4768
rect 7484 3738 7512 4762
rect 7576 4146 7604 4966
rect 7564 4140 7616 4146
rect 7564 4082 7616 4088
rect 7472 3732 7524 3738
rect 7472 3674 7524 3680
rect 6555 3292 6863 3301
rect 6555 3290 6561 3292
rect 6617 3290 6641 3292
rect 6697 3290 6721 3292
rect 6777 3290 6801 3292
rect 6857 3290 6863 3292
rect 6617 3238 6619 3290
rect 6799 3238 6801 3290
rect 6555 3236 6561 3238
rect 6617 3236 6641 3238
rect 6697 3236 6721 3238
rect 6777 3236 6801 3238
rect 6857 3236 6863 3238
rect 6555 3227 6863 3236
rect 6932 3194 6960 3454
rect 7288 3460 7340 3466
rect 7288 3402 7340 3408
rect 7012 3392 7064 3398
rect 7012 3334 7064 3340
rect 7024 3194 7052 3334
rect 7760 3210 7788 5102
rect 7873 4924 8181 4933
rect 7873 4922 7879 4924
rect 7935 4922 7959 4924
rect 8015 4922 8039 4924
rect 8095 4922 8119 4924
rect 8175 4922 8181 4924
rect 7935 4870 7937 4922
rect 8117 4870 8119 4922
rect 7873 4868 7879 4870
rect 7935 4868 7959 4870
rect 8015 4868 8039 4870
rect 8095 4868 8119 4870
rect 8175 4868 8181 4870
rect 7873 4859 8181 4868
rect 8220 4826 8248 5170
rect 8208 4820 8260 4826
rect 8208 4762 8260 4768
rect 8300 4616 8352 4622
rect 8300 4558 8352 4564
rect 8312 4078 8340 4558
rect 8404 4282 8432 5170
rect 8574 4584 8630 4593
rect 8574 4519 8576 4528
rect 8628 4519 8630 4528
rect 8576 4490 8628 4496
rect 8533 4380 8841 4389
rect 8533 4378 8539 4380
rect 8595 4378 8619 4380
rect 8675 4378 8699 4380
rect 8755 4378 8779 4380
rect 8835 4378 8841 4380
rect 8595 4326 8597 4378
rect 8777 4326 8779 4378
rect 8533 4324 8539 4326
rect 8595 4324 8619 4326
rect 8675 4324 8699 4326
rect 8755 4324 8779 4326
rect 8835 4324 8841 4326
rect 8533 4315 8841 4324
rect 8392 4276 8444 4282
rect 8392 4218 8444 4224
rect 8956 4146 8984 6054
rect 8944 4140 8996 4146
rect 8944 4082 8996 4088
rect 8300 4072 8352 4078
rect 8300 4014 8352 4020
rect 7873 3836 8181 3845
rect 7873 3834 7879 3836
rect 7935 3834 7959 3836
rect 8015 3834 8039 3836
rect 8095 3834 8119 3836
rect 8175 3834 8181 3836
rect 7935 3782 7937 3834
rect 8117 3782 8119 3834
rect 7873 3780 7879 3782
rect 7935 3780 7959 3782
rect 8015 3780 8039 3782
rect 8095 3780 8119 3782
rect 8175 3780 8181 3782
rect 7873 3771 8181 3780
rect 8022 3496 8078 3505
rect 8022 3431 8078 3440
rect 6736 3188 6788 3194
rect 6736 3130 6788 3136
rect 6920 3188 6972 3194
rect 6920 3130 6972 3136
rect 7012 3188 7064 3194
rect 7012 3130 7064 3136
rect 7392 3182 7788 3210
rect 8036 3194 8064 3431
rect 8312 3194 8340 4014
rect 8533 3292 8841 3301
rect 8533 3290 8539 3292
rect 8595 3290 8619 3292
rect 8675 3290 8699 3292
rect 8755 3290 8779 3292
rect 8835 3290 8841 3292
rect 8595 3238 8597 3290
rect 8777 3238 8779 3290
rect 8533 3236 8539 3238
rect 8595 3236 8619 3238
rect 8675 3236 8699 3238
rect 8755 3236 8779 3238
rect 8835 3236 8841 3238
rect 8533 3227 8841 3236
rect 8024 3188 8076 3194
rect 6460 2576 6512 2582
rect 6460 2518 6512 2524
rect 6368 2508 6420 2514
rect 6368 2450 6420 2456
rect 6748 2446 6776 3130
rect 7392 3126 7420 3182
rect 7380 3120 7432 3126
rect 6918 3088 6974 3097
rect 7380 3062 7432 3068
rect 6918 3023 6920 3032
rect 6972 3023 6974 3032
rect 7196 3052 7248 3058
rect 6920 2994 6972 3000
rect 7196 2994 7248 3000
rect 7012 2916 7064 2922
rect 7012 2858 7064 2864
rect 6828 2848 6880 2854
rect 6828 2790 6880 2796
rect 6840 2582 6868 2790
rect 7024 2650 7052 2858
rect 7012 2644 7064 2650
rect 7012 2586 7064 2592
rect 6828 2576 6880 2582
rect 6828 2518 6880 2524
rect 7208 2446 7236 2994
rect 7668 2854 7696 3182
rect 8024 3130 8076 3136
rect 8300 3188 8352 3194
rect 8300 3130 8352 3136
rect 7748 3052 7800 3058
rect 7748 2994 7800 3000
rect 7656 2848 7708 2854
rect 7656 2790 7708 2796
rect 7668 2582 7696 2790
rect 7656 2576 7708 2582
rect 7656 2518 7708 2524
rect 7760 2530 7788 2994
rect 8484 2984 8536 2990
rect 8390 2952 8446 2961
rect 8484 2926 8536 2932
rect 8390 2887 8446 2896
rect 8300 2848 8352 2854
rect 8300 2790 8352 2796
rect 7873 2748 8181 2757
rect 7873 2746 7879 2748
rect 7935 2746 7959 2748
rect 8015 2746 8039 2748
rect 8095 2746 8119 2748
rect 8175 2746 8181 2748
rect 7935 2694 7937 2746
rect 8117 2694 8119 2746
rect 7873 2692 7879 2694
rect 7935 2692 7959 2694
rect 8015 2692 8039 2694
rect 8095 2692 8119 2694
rect 8175 2692 8181 2694
rect 7873 2683 8181 2692
rect 8312 2582 8340 2790
rect 8300 2576 8352 2582
rect 7760 2502 7972 2530
rect 8300 2518 8352 2524
rect 7944 2446 7972 2502
rect 5816 2440 5868 2446
rect 5816 2382 5868 2388
rect 5908 2440 5960 2446
rect 5908 2382 5960 2388
rect 6736 2440 6788 2446
rect 6736 2382 6788 2388
rect 7196 2440 7248 2446
rect 7196 2382 7248 2388
rect 7932 2440 7984 2446
rect 7932 2382 7984 2388
rect 6460 2304 6512 2310
rect 6460 2246 6512 2252
rect 7472 2304 7524 2310
rect 7472 2246 7524 2252
rect 8024 2304 8076 2310
rect 8024 2246 8076 2252
rect 5356 2032 5408 2038
rect 5356 1974 5408 1980
rect 5724 2032 5776 2038
rect 5724 1974 5776 1980
rect 6472 1902 6500 2246
rect 6555 2204 6863 2213
rect 6555 2202 6561 2204
rect 6617 2202 6641 2204
rect 6697 2202 6721 2204
rect 6777 2202 6801 2204
rect 6857 2202 6863 2204
rect 6617 2150 6619 2202
rect 6799 2150 6801 2202
rect 6555 2148 6561 2150
rect 6617 2148 6641 2150
rect 6697 2148 6721 2150
rect 6777 2148 6801 2150
rect 6857 2148 6863 2150
rect 6555 2139 6863 2148
rect 3792 1896 3844 1902
rect 3792 1838 3844 1844
rect 6460 1896 6512 1902
rect 6460 1838 6512 1844
rect 7484 1766 7512 2246
rect 8036 2106 8064 2246
rect 8024 2100 8076 2106
rect 8024 2042 8076 2048
rect 3700 1760 3752 1766
rect 3700 1702 3752 1708
rect 7472 1760 7524 1766
rect 7472 1702 7524 1708
rect 8404 800 8432 2887
rect 8496 2582 8524 2926
rect 8484 2576 8536 2582
rect 8484 2518 8536 2524
rect 8533 2204 8841 2213
rect 8533 2202 8539 2204
rect 8595 2202 8619 2204
rect 8675 2202 8699 2204
rect 8755 2202 8779 2204
rect 8835 2202 8841 2204
rect 8595 2150 8597 2202
rect 8777 2150 8779 2202
rect 8533 2148 8539 2150
rect 8595 2148 8619 2150
rect 8675 2148 8699 2150
rect 8755 2148 8779 2150
rect 8835 2148 8841 2150
rect 8533 2139 8841 2148
rect 18 0 74 800
rect 8390 0 8446 800
<< via2 >>
rect 2605 9818 2661 9820
rect 2685 9818 2741 9820
rect 2765 9818 2821 9820
rect 2845 9818 2901 9820
rect 2605 9766 2651 9818
rect 2651 9766 2661 9818
rect 2685 9766 2715 9818
rect 2715 9766 2727 9818
rect 2727 9766 2741 9818
rect 2765 9766 2779 9818
rect 2779 9766 2791 9818
rect 2791 9766 2821 9818
rect 2845 9766 2855 9818
rect 2855 9766 2901 9818
rect 2605 9764 2661 9766
rect 2685 9764 2741 9766
rect 2765 9764 2821 9766
rect 2845 9764 2901 9766
rect 4583 9818 4639 9820
rect 4663 9818 4719 9820
rect 4743 9818 4799 9820
rect 4823 9818 4879 9820
rect 4583 9766 4629 9818
rect 4629 9766 4639 9818
rect 4663 9766 4693 9818
rect 4693 9766 4705 9818
rect 4705 9766 4719 9818
rect 4743 9766 4757 9818
rect 4757 9766 4769 9818
rect 4769 9766 4799 9818
rect 4823 9766 4833 9818
rect 4833 9766 4879 9818
rect 4583 9764 4639 9766
rect 4663 9764 4719 9766
rect 4743 9764 4799 9766
rect 4823 9764 4879 9766
rect 1945 9274 2001 9276
rect 2025 9274 2081 9276
rect 2105 9274 2161 9276
rect 2185 9274 2241 9276
rect 1945 9222 1991 9274
rect 1991 9222 2001 9274
rect 2025 9222 2055 9274
rect 2055 9222 2067 9274
rect 2067 9222 2081 9274
rect 2105 9222 2119 9274
rect 2119 9222 2131 9274
rect 2131 9222 2161 9274
rect 2185 9222 2195 9274
rect 2195 9222 2241 9274
rect 1945 9220 2001 9222
rect 2025 9220 2081 9222
rect 2105 9220 2161 9222
rect 2185 9220 2241 9222
rect 6561 9818 6617 9820
rect 6641 9818 6697 9820
rect 6721 9818 6777 9820
rect 6801 9818 6857 9820
rect 6561 9766 6607 9818
rect 6607 9766 6617 9818
rect 6641 9766 6671 9818
rect 6671 9766 6683 9818
rect 6683 9766 6697 9818
rect 6721 9766 6735 9818
rect 6735 9766 6747 9818
rect 6747 9766 6777 9818
rect 6801 9766 6811 9818
rect 6811 9766 6857 9818
rect 6561 9764 6617 9766
rect 6641 9764 6697 9766
rect 6721 9764 6777 9766
rect 6801 9764 6857 9766
rect 8539 9818 8595 9820
rect 8619 9818 8675 9820
rect 8699 9818 8755 9820
rect 8779 9818 8835 9820
rect 8539 9766 8585 9818
rect 8585 9766 8595 9818
rect 8619 9766 8649 9818
rect 8649 9766 8661 9818
rect 8661 9766 8675 9818
rect 8699 9766 8713 9818
rect 8713 9766 8725 9818
rect 8725 9766 8755 9818
rect 8779 9766 8789 9818
rect 8789 9766 8835 9818
rect 8539 9764 8595 9766
rect 8619 9764 8675 9766
rect 8699 9764 8755 9766
rect 8779 9764 8835 9766
rect 2605 8730 2661 8732
rect 2685 8730 2741 8732
rect 2765 8730 2821 8732
rect 2845 8730 2901 8732
rect 2605 8678 2651 8730
rect 2651 8678 2661 8730
rect 2685 8678 2715 8730
rect 2715 8678 2727 8730
rect 2727 8678 2741 8730
rect 2765 8678 2779 8730
rect 2779 8678 2791 8730
rect 2791 8678 2821 8730
rect 2845 8678 2855 8730
rect 2855 8678 2901 8730
rect 2605 8676 2661 8678
rect 2685 8676 2741 8678
rect 2765 8676 2821 8678
rect 2845 8676 2901 8678
rect 1945 8186 2001 8188
rect 2025 8186 2081 8188
rect 2105 8186 2161 8188
rect 2185 8186 2241 8188
rect 1945 8134 1991 8186
rect 1991 8134 2001 8186
rect 2025 8134 2055 8186
rect 2055 8134 2067 8186
rect 2067 8134 2081 8186
rect 2105 8134 2119 8186
rect 2119 8134 2131 8186
rect 2131 8134 2161 8186
rect 2185 8134 2195 8186
rect 2195 8134 2241 8186
rect 1945 8132 2001 8134
rect 2025 8132 2081 8134
rect 2105 8132 2161 8134
rect 2185 8132 2241 8134
rect 1945 7098 2001 7100
rect 2025 7098 2081 7100
rect 2105 7098 2161 7100
rect 2185 7098 2241 7100
rect 1945 7046 1991 7098
rect 1991 7046 2001 7098
rect 2025 7046 2055 7098
rect 2055 7046 2067 7098
rect 2067 7046 2081 7098
rect 2105 7046 2119 7098
rect 2119 7046 2131 7098
rect 2131 7046 2161 7098
rect 2185 7046 2195 7098
rect 2195 7046 2241 7098
rect 1945 7044 2001 7046
rect 2025 7044 2081 7046
rect 2105 7044 2161 7046
rect 2185 7044 2241 7046
rect 1766 6316 1822 6352
rect 1766 6296 1768 6316
rect 1768 6296 1820 6316
rect 1820 6296 1822 6316
rect 2605 7642 2661 7644
rect 2685 7642 2741 7644
rect 2765 7642 2821 7644
rect 2845 7642 2901 7644
rect 2605 7590 2651 7642
rect 2651 7590 2661 7642
rect 2685 7590 2715 7642
rect 2715 7590 2727 7642
rect 2727 7590 2741 7642
rect 2765 7590 2779 7642
rect 2779 7590 2791 7642
rect 2791 7590 2821 7642
rect 2845 7590 2855 7642
rect 2855 7590 2901 7642
rect 2605 7588 2661 7590
rect 2685 7588 2741 7590
rect 2765 7588 2821 7590
rect 2845 7588 2901 7590
rect 2605 6554 2661 6556
rect 2685 6554 2741 6556
rect 2765 6554 2821 6556
rect 2845 6554 2901 6556
rect 2605 6502 2651 6554
rect 2651 6502 2661 6554
rect 2685 6502 2715 6554
rect 2715 6502 2727 6554
rect 2727 6502 2741 6554
rect 2765 6502 2779 6554
rect 2779 6502 2791 6554
rect 2791 6502 2821 6554
rect 2845 6502 2855 6554
rect 2855 6502 2901 6554
rect 2605 6500 2661 6502
rect 2685 6500 2741 6502
rect 2765 6500 2821 6502
rect 2845 6500 2901 6502
rect 3606 8880 3662 8936
rect 1945 6010 2001 6012
rect 2025 6010 2081 6012
rect 2105 6010 2161 6012
rect 2185 6010 2241 6012
rect 1945 5958 1991 6010
rect 1991 5958 2001 6010
rect 2025 5958 2055 6010
rect 2055 5958 2067 6010
rect 2067 5958 2081 6010
rect 2105 5958 2119 6010
rect 2119 5958 2131 6010
rect 2131 5958 2161 6010
rect 2185 5958 2195 6010
rect 2195 5958 2241 6010
rect 1945 5956 2001 5958
rect 2025 5956 2081 5958
rect 2105 5956 2161 5958
rect 2185 5956 2241 5958
rect 2870 6160 2926 6216
rect 1945 4922 2001 4924
rect 2025 4922 2081 4924
rect 2105 4922 2161 4924
rect 2185 4922 2241 4924
rect 1945 4870 1991 4922
rect 1991 4870 2001 4922
rect 2025 4870 2055 4922
rect 2055 4870 2067 4922
rect 2067 4870 2081 4922
rect 2105 4870 2119 4922
rect 2119 4870 2131 4922
rect 2131 4870 2161 4922
rect 2185 4870 2195 4922
rect 2195 4870 2241 4922
rect 1945 4868 2001 4870
rect 2025 4868 2081 4870
rect 2105 4868 2161 4870
rect 2185 4868 2241 4870
rect 2134 4664 2190 4720
rect 2605 5466 2661 5468
rect 2685 5466 2741 5468
rect 2765 5466 2821 5468
rect 2845 5466 2901 5468
rect 2605 5414 2651 5466
rect 2651 5414 2661 5466
rect 2685 5414 2715 5466
rect 2715 5414 2727 5466
rect 2727 5414 2741 5466
rect 2765 5414 2779 5466
rect 2779 5414 2791 5466
rect 2791 5414 2821 5466
rect 2845 5414 2855 5466
rect 2855 5414 2901 5466
rect 2605 5412 2661 5414
rect 2685 5412 2741 5414
rect 2765 5412 2821 5414
rect 2845 5412 2901 5414
rect 2870 4800 2926 4856
rect 2605 4378 2661 4380
rect 2685 4378 2741 4380
rect 2765 4378 2821 4380
rect 2845 4378 2901 4380
rect 2605 4326 2651 4378
rect 2651 4326 2661 4378
rect 2685 4326 2715 4378
rect 2715 4326 2727 4378
rect 2727 4326 2741 4378
rect 2765 4326 2779 4378
rect 2779 4326 2791 4378
rect 2791 4326 2821 4378
rect 2845 4326 2855 4378
rect 2855 4326 2901 4378
rect 2605 4324 2661 4326
rect 2685 4324 2741 4326
rect 2765 4324 2821 4326
rect 2845 4324 2901 4326
rect 1490 3440 1546 3496
rect 1766 4004 1822 4040
rect 1766 3984 1768 4004
rect 1768 3984 1820 4004
rect 1820 3984 1822 4004
rect 1945 3834 2001 3836
rect 2025 3834 2081 3836
rect 2105 3834 2161 3836
rect 2185 3834 2241 3836
rect 1945 3782 1991 3834
rect 1991 3782 2001 3834
rect 2025 3782 2055 3834
rect 2055 3782 2067 3834
rect 2067 3782 2081 3834
rect 2105 3782 2119 3834
rect 2119 3782 2131 3834
rect 2131 3782 2161 3834
rect 2185 3782 2195 3834
rect 2195 3782 2241 3834
rect 1945 3780 2001 3782
rect 2025 3780 2081 3782
rect 2105 3780 2161 3782
rect 2185 3780 2241 3782
rect 2042 2896 2098 2952
rect 3923 9274 3979 9276
rect 4003 9274 4059 9276
rect 4083 9274 4139 9276
rect 4163 9274 4219 9276
rect 3923 9222 3969 9274
rect 3969 9222 3979 9274
rect 4003 9222 4033 9274
rect 4033 9222 4045 9274
rect 4045 9222 4059 9274
rect 4083 9222 4097 9274
rect 4097 9222 4109 9274
rect 4109 9222 4139 9274
rect 4163 9222 4173 9274
rect 4173 9222 4219 9274
rect 3923 9220 3979 9222
rect 4003 9220 4059 9222
rect 4083 9220 4139 9222
rect 4163 9220 4219 9222
rect 3923 8186 3979 8188
rect 4003 8186 4059 8188
rect 4083 8186 4139 8188
rect 4163 8186 4219 8188
rect 3923 8134 3969 8186
rect 3969 8134 3979 8186
rect 4003 8134 4033 8186
rect 4033 8134 4045 8186
rect 4045 8134 4059 8186
rect 4083 8134 4097 8186
rect 4097 8134 4109 8186
rect 4109 8134 4139 8186
rect 4163 8134 4173 8186
rect 4173 8134 4219 8186
rect 3923 8132 3979 8134
rect 4003 8132 4059 8134
rect 4083 8132 4139 8134
rect 4163 8132 4219 8134
rect 4583 8730 4639 8732
rect 4663 8730 4719 8732
rect 4743 8730 4799 8732
rect 4823 8730 4879 8732
rect 4583 8678 4629 8730
rect 4629 8678 4639 8730
rect 4663 8678 4693 8730
rect 4693 8678 4705 8730
rect 4705 8678 4719 8730
rect 4743 8678 4757 8730
rect 4757 8678 4769 8730
rect 4769 8678 4799 8730
rect 4823 8678 4833 8730
rect 4833 8678 4879 8730
rect 4583 8676 4639 8678
rect 4663 8676 4719 8678
rect 4743 8676 4799 8678
rect 4823 8676 4879 8678
rect 3923 7098 3979 7100
rect 4003 7098 4059 7100
rect 4083 7098 4139 7100
rect 4163 7098 4219 7100
rect 3923 7046 3969 7098
rect 3969 7046 3979 7098
rect 4003 7046 4033 7098
rect 4033 7046 4045 7098
rect 4045 7046 4059 7098
rect 4083 7046 4097 7098
rect 4097 7046 4109 7098
rect 4109 7046 4139 7098
rect 4163 7046 4173 7098
rect 4173 7046 4219 7098
rect 3923 7044 3979 7046
rect 4003 7044 4059 7046
rect 4083 7044 4139 7046
rect 4163 7044 4219 7046
rect 3882 6160 3938 6216
rect 3923 6010 3979 6012
rect 4003 6010 4059 6012
rect 4083 6010 4139 6012
rect 4163 6010 4219 6012
rect 3923 5958 3969 6010
rect 3969 5958 3979 6010
rect 4003 5958 4033 6010
rect 4033 5958 4045 6010
rect 4045 5958 4059 6010
rect 4083 5958 4097 6010
rect 4097 5958 4109 6010
rect 4109 5958 4139 6010
rect 4163 5958 4173 6010
rect 4173 5958 4219 6010
rect 3923 5956 3979 5958
rect 4003 5956 4059 5958
rect 4083 5956 4139 5958
rect 4163 5956 4219 5958
rect 3882 5752 3938 5808
rect 4158 5652 4160 5672
rect 4160 5652 4212 5672
rect 4212 5652 4214 5672
rect 4158 5616 4214 5652
rect 3923 4922 3979 4924
rect 4003 4922 4059 4924
rect 4083 4922 4139 4924
rect 4163 4922 4219 4924
rect 3923 4870 3969 4922
rect 3969 4870 3979 4922
rect 4003 4870 4033 4922
rect 4033 4870 4045 4922
rect 4045 4870 4059 4922
rect 4083 4870 4097 4922
rect 4097 4870 4109 4922
rect 4109 4870 4139 4922
rect 4163 4870 4173 4922
rect 4173 4870 4219 4922
rect 3923 4868 3979 4870
rect 4003 4868 4059 4870
rect 4083 4868 4139 4870
rect 4163 4868 4219 4870
rect 4066 4564 4068 4584
rect 4068 4564 4120 4584
rect 4120 4564 4122 4584
rect 4066 4528 4122 4564
rect 2605 3290 2661 3292
rect 2685 3290 2741 3292
rect 2765 3290 2821 3292
rect 2845 3290 2901 3292
rect 2605 3238 2651 3290
rect 2651 3238 2661 3290
rect 2685 3238 2715 3290
rect 2715 3238 2727 3290
rect 2727 3238 2741 3290
rect 2765 3238 2779 3290
rect 2779 3238 2791 3290
rect 2791 3238 2821 3290
rect 2845 3238 2855 3290
rect 2855 3238 2901 3290
rect 2605 3236 2661 3238
rect 2685 3236 2741 3238
rect 2765 3236 2821 3238
rect 2845 3236 2901 3238
rect 1945 2746 2001 2748
rect 2025 2746 2081 2748
rect 2105 2746 2161 2748
rect 2185 2746 2241 2748
rect 1945 2694 1991 2746
rect 1991 2694 2001 2746
rect 2025 2694 2055 2746
rect 2055 2694 2067 2746
rect 2067 2694 2081 2746
rect 2105 2694 2119 2746
rect 2119 2694 2131 2746
rect 2131 2694 2161 2746
rect 2185 2694 2195 2746
rect 2195 2694 2241 2746
rect 1945 2692 2001 2694
rect 2025 2692 2081 2694
rect 2105 2692 2161 2694
rect 2185 2692 2241 2694
rect 3238 3032 3294 3088
rect 2502 2488 2558 2544
rect 3923 3834 3979 3836
rect 4003 3834 4059 3836
rect 4083 3834 4139 3836
rect 4163 3834 4219 3836
rect 3923 3782 3969 3834
rect 3969 3782 3979 3834
rect 4003 3782 4033 3834
rect 4033 3782 4045 3834
rect 4045 3782 4059 3834
rect 4083 3782 4097 3834
rect 4097 3782 4109 3834
rect 4109 3782 4139 3834
rect 4163 3782 4173 3834
rect 4173 3782 4219 3834
rect 3923 3780 3979 3782
rect 4003 3780 4059 3782
rect 4083 3780 4139 3782
rect 4163 3780 4219 3782
rect 3974 3576 4030 3632
rect 3422 2388 3424 2408
rect 3424 2388 3476 2408
rect 3476 2388 3478 2408
rect 3422 2352 3478 2388
rect 2605 2202 2661 2204
rect 2685 2202 2741 2204
rect 2765 2202 2821 2204
rect 2845 2202 2901 2204
rect 2605 2150 2651 2202
rect 2651 2150 2661 2202
rect 2685 2150 2715 2202
rect 2715 2150 2727 2202
rect 2727 2150 2741 2202
rect 2765 2150 2779 2202
rect 2779 2150 2791 2202
rect 2791 2150 2821 2202
rect 2845 2150 2855 2202
rect 2855 2150 2901 2202
rect 2605 2148 2661 2150
rect 2685 2148 2741 2150
rect 2765 2148 2821 2150
rect 2845 2148 2901 2150
rect 3923 2746 3979 2748
rect 4003 2746 4059 2748
rect 4083 2746 4139 2748
rect 4163 2746 4219 2748
rect 3923 2694 3969 2746
rect 3969 2694 3979 2746
rect 4003 2694 4033 2746
rect 4033 2694 4045 2746
rect 4045 2694 4059 2746
rect 4083 2694 4097 2746
rect 4097 2694 4109 2746
rect 4109 2694 4139 2746
rect 4163 2694 4173 2746
rect 4173 2694 4219 2746
rect 3923 2692 3979 2694
rect 4003 2692 4059 2694
rect 4083 2692 4139 2694
rect 4163 2692 4219 2694
rect 4583 7642 4639 7644
rect 4663 7642 4719 7644
rect 4743 7642 4799 7644
rect 4823 7642 4879 7644
rect 4583 7590 4629 7642
rect 4629 7590 4639 7642
rect 4663 7590 4693 7642
rect 4693 7590 4705 7642
rect 4705 7590 4719 7642
rect 4743 7590 4757 7642
rect 4757 7590 4769 7642
rect 4769 7590 4799 7642
rect 4823 7590 4833 7642
rect 4833 7590 4879 7642
rect 4583 7588 4639 7590
rect 4663 7588 4719 7590
rect 4743 7588 4799 7590
rect 4823 7588 4879 7590
rect 4583 6554 4639 6556
rect 4663 6554 4719 6556
rect 4743 6554 4799 6556
rect 4823 6554 4879 6556
rect 4583 6502 4629 6554
rect 4629 6502 4639 6554
rect 4663 6502 4693 6554
rect 4693 6502 4705 6554
rect 4705 6502 4719 6554
rect 4743 6502 4757 6554
rect 4757 6502 4769 6554
rect 4769 6502 4799 6554
rect 4823 6502 4833 6554
rect 4833 6502 4879 6554
rect 4583 6500 4639 6502
rect 4663 6500 4719 6502
rect 4743 6500 4799 6502
rect 4823 6500 4879 6502
rect 4526 6316 4582 6352
rect 4526 6296 4528 6316
rect 4528 6296 4580 6316
rect 4580 6296 4582 6316
rect 5078 7828 5080 7848
rect 5080 7828 5132 7848
rect 5132 7828 5134 7848
rect 5078 7792 5134 7828
rect 5901 9274 5957 9276
rect 5981 9274 6037 9276
rect 6061 9274 6117 9276
rect 6141 9274 6197 9276
rect 5901 9222 5947 9274
rect 5947 9222 5957 9274
rect 5981 9222 6011 9274
rect 6011 9222 6023 9274
rect 6023 9222 6037 9274
rect 6061 9222 6075 9274
rect 6075 9222 6087 9274
rect 6087 9222 6117 9274
rect 6141 9222 6151 9274
rect 6151 9222 6197 9274
rect 5901 9220 5957 9222
rect 5981 9220 6037 9222
rect 6061 9220 6117 9222
rect 6141 9220 6197 9222
rect 5170 5888 5226 5944
rect 4583 5466 4639 5468
rect 4663 5466 4719 5468
rect 4743 5466 4799 5468
rect 4823 5466 4879 5468
rect 4583 5414 4629 5466
rect 4629 5414 4639 5466
rect 4663 5414 4693 5466
rect 4693 5414 4705 5466
rect 4705 5414 4719 5466
rect 4743 5414 4757 5466
rect 4757 5414 4769 5466
rect 4769 5414 4799 5466
rect 4823 5414 4833 5466
rect 4833 5414 4879 5466
rect 4583 5412 4639 5414
rect 4663 5412 4719 5414
rect 4743 5412 4799 5414
rect 4823 5412 4879 5414
rect 4618 4800 4674 4856
rect 4802 4664 4858 4720
rect 4986 5344 5042 5400
rect 5170 5072 5226 5128
rect 4583 4378 4639 4380
rect 4663 4378 4719 4380
rect 4743 4378 4799 4380
rect 4823 4378 4879 4380
rect 4583 4326 4629 4378
rect 4629 4326 4639 4378
rect 4663 4326 4693 4378
rect 4693 4326 4705 4378
rect 4705 4326 4719 4378
rect 4743 4326 4757 4378
rect 4757 4326 4769 4378
rect 4769 4326 4799 4378
rect 4823 4326 4833 4378
rect 4833 4326 4879 4378
rect 4583 4324 4639 4326
rect 4663 4324 4719 4326
rect 4743 4324 4799 4326
rect 4823 4324 4879 4326
rect 5078 4936 5134 4992
rect 5901 8186 5957 8188
rect 5981 8186 6037 8188
rect 6061 8186 6117 8188
rect 6141 8186 6197 8188
rect 5901 8134 5947 8186
rect 5947 8134 5957 8186
rect 5981 8134 6011 8186
rect 6011 8134 6023 8186
rect 6023 8134 6037 8186
rect 6061 8134 6075 8186
rect 6075 8134 6087 8186
rect 6087 8134 6117 8186
rect 6141 8134 6151 8186
rect 6151 8134 6197 8186
rect 5901 8132 5957 8134
rect 5981 8132 6037 8134
rect 6061 8132 6117 8134
rect 6141 8132 6197 8134
rect 5906 7928 5962 7984
rect 5630 7248 5686 7304
rect 6090 7248 6146 7304
rect 6366 8336 6422 8392
rect 6366 7792 6422 7848
rect 6561 8730 6617 8732
rect 6641 8730 6697 8732
rect 6721 8730 6777 8732
rect 6801 8730 6857 8732
rect 6561 8678 6607 8730
rect 6607 8678 6617 8730
rect 6641 8678 6671 8730
rect 6671 8678 6683 8730
rect 6683 8678 6697 8730
rect 6721 8678 6735 8730
rect 6735 8678 6747 8730
rect 6747 8678 6777 8730
rect 6801 8678 6811 8730
rect 6811 8678 6857 8730
rect 6561 8676 6617 8678
rect 6641 8676 6697 8678
rect 6721 8676 6777 8678
rect 6801 8676 6857 8678
rect 6561 7642 6617 7644
rect 6641 7642 6697 7644
rect 6721 7642 6777 7644
rect 6801 7642 6857 7644
rect 6561 7590 6607 7642
rect 6607 7590 6617 7642
rect 6641 7590 6671 7642
rect 6671 7590 6683 7642
rect 6683 7590 6697 7642
rect 6721 7590 6735 7642
rect 6735 7590 6747 7642
rect 6747 7590 6777 7642
rect 6801 7590 6811 7642
rect 6811 7590 6857 7642
rect 6561 7588 6617 7590
rect 6641 7588 6697 7590
rect 6721 7588 6777 7590
rect 6801 7588 6857 7590
rect 5901 7098 5957 7100
rect 5981 7098 6037 7100
rect 6061 7098 6117 7100
rect 6141 7098 6197 7100
rect 5901 7046 5947 7098
rect 5947 7046 5957 7098
rect 5981 7046 6011 7098
rect 6011 7046 6023 7098
rect 6023 7046 6037 7098
rect 6061 7046 6075 7098
rect 6075 7046 6087 7098
rect 6087 7046 6117 7098
rect 6141 7046 6151 7098
rect 6151 7046 6197 7098
rect 5901 7044 5957 7046
rect 5981 7044 6037 7046
rect 6061 7044 6117 7046
rect 6141 7044 6197 7046
rect 5901 6010 5957 6012
rect 5981 6010 6037 6012
rect 6061 6010 6117 6012
rect 6141 6010 6197 6012
rect 5901 5958 5947 6010
rect 5947 5958 5957 6010
rect 5981 5958 6011 6010
rect 6011 5958 6023 6010
rect 6023 5958 6037 6010
rect 6061 5958 6075 6010
rect 6075 5958 6087 6010
rect 6087 5958 6117 6010
rect 6141 5958 6151 6010
rect 6151 5958 6197 6010
rect 5901 5956 5957 5958
rect 5981 5956 6037 5958
rect 6061 5956 6117 5958
rect 6141 5956 6197 5958
rect 5538 5616 5594 5672
rect 5262 4800 5318 4856
rect 5262 4392 5318 4448
rect 5170 3612 5172 3632
rect 5172 3612 5224 3632
rect 5224 3612 5226 3632
rect 5170 3576 5226 3612
rect 4583 3290 4639 3292
rect 4663 3290 4719 3292
rect 4743 3290 4799 3292
rect 4823 3290 4879 3292
rect 4583 3238 4629 3290
rect 4629 3238 4639 3290
rect 4663 3238 4693 3290
rect 4693 3238 4705 3290
rect 4705 3238 4719 3290
rect 4743 3238 4757 3290
rect 4757 3238 4769 3290
rect 4769 3238 4799 3290
rect 4823 3238 4833 3290
rect 4833 3238 4879 3290
rect 4583 3236 4639 3238
rect 4663 3236 4719 3238
rect 4743 3236 4799 3238
rect 4823 3236 4879 3238
rect 5078 2488 5134 2544
rect 4583 2202 4639 2204
rect 4663 2202 4719 2204
rect 4743 2202 4799 2204
rect 4823 2202 4879 2204
rect 4583 2150 4629 2202
rect 4629 2150 4639 2202
rect 4663 2150 4693 2202
rect 4693 2150 4705 2202
rect 4705 2150 4719 2202
rect 4743 2150 4757 2202
rect 4757 2150 4769 2202
rect 4769 2150 4799 2202
rect 4823 2150 4833 2202
rect 4833 2150 4879 2202
rect 4583 2148 4639 2150
rect 4663 2148 4719 2150
rect 4743 2148 4799 2150
rect 4823 2148 4879 2150
rect 5630 4936 5686 4992
rect 5630 2388 5632 2408
rect 5632 2388 5684 2408
rect 5684 2388 5686 2408
rect 5630 2352 5686 2388
rect 7879 9274 7935 9276
rect 7959 9274 8015 9276
rect 8039 9274 8095 9276
rect 8119 9274 8175 9276
rect 7879 9222 7925 9274
rect 7925 9222 7935 9274
rect 7959 9222 7989 9274
rect 7989 9222 8001 9274
rect 8001 9222 8015 9274
rect 8039 9222 8053 9274
rect 8053 9222 8065 9274
rect 8065 9222 8095 9274
rect 8119 9222 8129 9274
rect 8129 9222 8175 9274
rect 7879 9220 7935 9222
rect 7959 9220 8015 9222
rect 8039 9220 8095 9222
rect 8119 9220 8175 9222
rect 6561 6554 6617 6556
rect 6641 6554 6697 6556
rect 6721 6554 6777 6556
rect 6801 6554 6857 6556
rect 6561 6502 6607 6554
rect 6607 6502 6617 6554
rect 6641 6502 6671 6554
rect 6671 6502 6683 6554
rect 6683 6502 6697 6554
rect 6721 6502 6735 6554
rect 6735 6502 6747 6554
rect 6747 6502 6777 6554
rect 6801 6502 6811 6554
rect 6811 6502 6857 6554
rect 6561 6500 6617 6502
rect 6641 6500 6697 6502
rect 6721 6500 6777 6502
rect 6801 6500 6857 6502
rect 6090 5072 6146 5128
rect 5901 4922 5957 4924
rect 5981 4922 6037 4924
rect 6061 4922 6117 4924
rect 6141 4922 6197 4924
rect 5901 4870 5947 4922
rect 5947 4870 5957 4922
rect 5981 4870 6011 4922
rect 6011 4870 6023 4922
rect 6023 4870 6037 4922
rect 6061 4870 6075 4922
rect 6075 4870 6087 4922
rect 6087 4870 6117 4922
rect 6141 4870 6151 4922
rect 6151 4870 6197 4922
rect 5901 4868 5957 4870
rect 5981 4868 6037 4870
rect 6061 4868 6117 4870
rect 6141 4868 6197 4870
rect 5998 4528 6054 4584
rect 5901 3834 5957 3836
rect 5981 3834 6037 3836
rect 6061 3834 6117 3836
rect 6141 3834 6197 3836
rect 5901 3782 5947 3834
rect 5947 3782 5957 3834
rect 5981 3782 6011 3834
rect 6011 3782 6023 3834
rect 6023 3782 6037 3834
rect 6061 3782 6075 3834
rect 6075 3782 6087 3834
rect 6087 3782 6117 3834
rect 6141 3782 6151 3834
rect 6151 3782 6197 3834
rect 5901 3780 5957 3782
rect 5981 3780 6037 3782
rect 6061 3780 6117 3782
rect 6141 3780 6197 3782
rect 6561 5466 6617 5468
rect 6641 5466 6697 5468
rect 6721 5466 6777 5468
rect 6801 5466 6857 5468
rect 6561 5414 6607 5466
rect 6607 5414 6617 5466
rect 6641 5414 6671 5466
rect 6671 5414 6683 5466
rect 6683 5414 6697 5466
rect 6721 5414 6735 5466
rect 6735 5414 6747 5466
rect 6747 5414 6777 5466
rect 6801 5414 6811 5466
rect 6811 5414 6857 5466
rect 6561 5412 6617 5414
rect 6641 5412 6697 5414
rect 6721 5412 6777 5414
rect 6801 5412 6857 5414
rect 6458 5208 6514 5264
rect 6642 5092 6698 5128
rect 6642 5072 6644 5092
rect 6644 5072 6696 5092
rect 6696 5072 6698 5092
rect 8539 8730 8595 8732
rect 8619 8730 8675 8732
rect 8699 8730 8755 8732
rect 8779 8730 8835 8732
rect 8539 8678 8585 8730
rect 8585 8678 8595 8730
rect 8619 8678 8649 8730
rect 8649 8678 8661 8730
rect 8661 8678 8675 8730
rect 8699 8678 8713 8730
rect 8713 8678 8725 8730
rect 8725 8678 8755 8730
rect 8779 8678 8789 8730
rect 8789 8678 8835 8730
rect 8539 8676 8595 8678
rect 8619 8676 8675 8678
rect 8699 8676 8755 8678
rect 8779 8676 8835 8678
rect 7879 8186 7935 8188
rect 7959 8186 8015 8188
rect 8039 8186 8095 8188
rect 8119 8186 8175 8188
rect 7879 8134 7925 8186
rect 7925 8134 7935 8186
rect 7959 8134 7989 8186
rect 7989 8134 8001 8186
rect 8001 8134 8015 8186
rect 8039 8134 8053 8186
rect 8053 8134 8065 8186
rect 8065 8134 8095 8186
rect 8119 8134 8129 8186
rect 8129 8134 8175 8186
rect 7879 8132 7935 8134
rect 7959 8132 8015 8134
rect 8039 8132 8095 8134
rect 8119 8132 8175 8134
rect 7562 7948 7618 7984
rect 7562 7928 7564 7948
rect 7564 7928 7616 7948
rect 7616 7928 7618 7948
rect 8114 7928 8170 7984
rect 6458 4664 6514 4720
rect 6561 4378 6617 4380
rect 6641 4378 6697 4380
rect 6721 4378 6777 4380
rect 6801 4378 6857 4380
rect 6561 4326 6607 4378
rect 6607 4326 6617 4378
rect 6641 4326 6671 4378
rect 6671 4326 6683 4378
rect 6683 4326 6697 4378
rect 6721 4326 6735 4378
rect 6735 4326 6747 4378
rect 6747 4326 6777 4378
rect 6801 4326 6811 4378
rect 6811 4326 6857 4378
rect 6561 4324 6617 4326
rect 6641 4324 6697 4326
rect 6721 4324 6777 4326
rect 6801 4324 6857 4326
rect 7010 4256 7066 4312
rect 5901 2746 5957 2748
rect 5981 2746 6037 2748
rect 6061 2746 6117 2748
rect 6141 2746 6197 2748
rect 5901 2694 5947 2746
rect 5947 2694 5957 2746
rect 5981 2694 6011 2746
rect 6011 2694 6023 2746
rect 6023 2694 6037 2746
rect 6061 2694 6075 2746
rect 6075 2694 6087 2746
rect 6087 2694 6117 2746
rect 6141 2694 6151 2746
rect 6151 2694 6197 2746
rect 5901 2692 5957 2694
rect 5981 2692 6037 2694
rect 6061 2692 6117 2694
rect 6141 2692 6197 2694
rect 7879 7098 7935 7100
rect 7959 7098 8015 7100
rect 8039 7098 8095 7100
rect 8119 7098 8175 7100
rect 7879 7046 7925 7098
rect 7925 7046 7935 7098
rect 7959 7046 7989 7098
rect 7989 7046 8001 7098
rect 8001 7046 8015 7098
rect 8039 7046 8053 7098
rect 8053 7046 8065 7098
rect 8065 7046 8095 7098
rect 8119 7046 8129 7098
rect 8129 7046 8175 7098
rect 7879 7044 7935 7046
rect 7959 7044 8015 7046
rect 8039 7044 8095 7046
rect 8119 7044 8175 7046
rect 8539 7642 8595 7644
rect 8619 7642 8675 7644
rect 8699 7642 8755 7644
rect 8779 7642 8835 7644
rect 8539 7590 8585 7642
rect 8585 7590 8595 7642
rect 8619 7590 8649 7642
rect 8649 7590 8661 7642
rect 8661 7590 8675 7642
rect 8699 7590 8713 7642
rect 8713 7590 8725 7642
rect 8725 7590 8755 7642
rect 8779 7590 8789 7642
rect 8789 7590 8835 7642
rect 8539 7588 8595 7590
rect 8619 7588 8675 7590
rect 8699 7588 8755 7590
rect 8779 7588 8835 7590
rect 9034 7520 9090 7576
rect 7879 6010 7935 6012
rect 7959 6010 8015 6012
rect 8039 6010 8095 6012
rect 8119 6010 8175 6012
rect 7879 5958 7925 6010
rect 7925 5958 7935 6010
rect 7959 5958 7989 6010
rect 7989 5958 8001 6010
rect 8001 5958 8015 6010
rect 8039 5958 8053 6010
rect 8053 5958 8065 6010
rect 8065 5958 8095 6010
rect 8119 5958 8129 6010
rect 8129 5958 8175 6010
rect 7879 5956 7935 5958
rect 7959 5956 8015 5958
rect 8039 5956 8095 5958
rect 8119 5956 8175 5958
rect 8539 6554 8595 6556
rect 8619 6554 8675 6556
rect 8699 6554 8755 6556
rect 8779 6554 8835 6556
rect 8539 6502 8585 6554
rect 8585 6502 8595 6554
rect 8619 6502 8649 6554
rect 8649 6502 8661 6554
rect 8661 6502 8675 6554
rect 8699 6502 8713 6554
rect 8713 6502 8725 6554
rect 8725 6502 8755 6554
rect 8779 6502 8789 6554
rect 8789 6502 8835 6554
rect 8539 6500 8595 6502
rect 8619 6500 8675 6502
rect 8699 6500 8755 6502
rect 8779 6500 8835 6502
rect 8539 5466 8595 5468
rect 8619 5466 8675 5468
rect 8699 5466 8755 5468
rect 8779 5466 8835 5468
rect 8539 5414 8585 5466
rect 8585 5414 8595 5466
rect 8619 5414 8649 5466
rect 8649 5414 8661 5466
rect 8661 5414 8675 5466
rect 8699 5414 8713 5466
rect 8713 5414 8725 5466
rect 8725 5414 8755 5466
rect 8779 5414 8789 5466
rect 8789 5414 8835 5466
rect 8539 5412 8595 5414
rect 8619 5412 8675 5414
rect 8699 5412 8755 5414
rect 8779 5412 8835 5414
rect 6561 3290 6617 3292
rect 6641 3290 6697 3292
rect 6721 3290 6777 3292
rect 6801 3290 6857 3292
rect 6561 3238 6607 3290
rect 6607 3238 6617 3290
rect 6641 3238 6671 3290
rect 6671 3238 6683 3290
rect 6683 3238 6697 3290
rect 6721 3238 6735 3290
rect 6735 3238 6747 3290
rect 6747 3238 6777 3290
rect 6801 3238 6811 3290
rect 6811 3238 6857 3290
rect 6561 3236 6617 3238
rect 6641 3236 6697 3238
rect 6721 3236 6777 3238
rect 6801 3236 6857 3238
rect 7879 4922 7935 4924
rect 7959 4922 8015 4924
rect 8039 4922 8095 4924
rect 8119 4922 8175 4924
rect 7879 4870 7925 4922
rect 7925 4870 7935 4922
rect 7959 4870 7989 4922
rect 7989 4870 8001 4922
rect 8001 4870 8015 4922
rect 8039 4870 8053 4922
rect 8053 4870 8065 4922
rect 8065 4870 8095 4922
rect 8119 4870 8129 4922
rect 8129 4870 8175 4922
rect 7879 4868 7935 4870
rect 7959 4868 8015 4870
rect 8039 4868 8095 4870
rect 8119 4868 8175 4870
rect 8574 4548 8630 4584
rect 8574 4528 8576 4548
rect 8576 4528 8628 4548
rect 8628 4528 8630 4548
rect 8539 4378 8595 4380
rect 8619 4378 8675 4380
rect 8699 4378 8755 4380
rect 8779 4378 8835 4380
rect 8539 4326 8585 4378
rect 8585 4326 8595 4378
rect 8619 4326 8649 4378
rect 8649 4326 8661 4378
rect 8661 4326 8675 4378
rect 8699 4326 8713 4378
rect 8713 4326 8725 4378
rect 8725 4326 8755 4378
rect 8779 4326 8789 4378
rect 8789 4326 8835 4378
rect 8539 4324 8595 4326
rect 8619 4324 8675 4326
rect 8699 4324 8755 4326
rect 8779 4324 8835 4326
rect 7879 3834 7935 3836
rect 7959 3834 8015 3836
rect 8039 3834 8095 3836
rect 8119 3834 8175 3836
rect 7879 3782 7925 3834
rect 7925 3782 7935 3834
rect 7959 3782 7989 3834
rect 7989 3782 8001 3834
rect 8001 3782 8015 3834
rect 8039 3782 8053 3834
rect 8053 3782 8065 3834
rect 8065 3782 8095 3834
rect 8119 3782 8129 3834
rect 8129 3782 8175 3834
rect 7879 3780 7935 3782
rect 7959 3780 8015 3782
rect 8039 3780 8095 3782
rect 8119 3780 8175 3782
rect 8022 3440 8078 3496
rect 8539 3290 8595 3292
rect 8619 3290 8675 3292
rect 8699 3290 8755 3292
rect 8779 3290 8835 3292
rect 8539 3238 8585 3290
rect 8585 3238 8595 3290
rect 8619 3238 8649 3290
rect 8649 3238 8661 3290
rect 8661 3238 8675 3290
rect 8699 3238 8713 3290
rect 8713 3238 8725 3290
rect 8725 3238 8755 3290
rect 8779 3238 8789 3290
rect 8789 3238 8835 3290
rect 8539 3236 8595 3238
rect 8619 3236 8675 3238
rect 8699 3236 8755 3238
rect 8779 3236 8835 3238
rect 6918 3052 6974 3088
rect 6918 3032 6920 3052
rect 6920 3032 6972 3052
rect 6972 3032 6974 3052
rect 8390 2896 8446 2952
rect 7879 2746 7935 2748
rect 7959 2746 8015 2748
rect 8039 2746 8095 2748
rect 8119 2746 8175 2748
rect 7879 2694 7925 2746
rect 7925 2694 7935 2746
rect 7959 2694 7989 2746
rect 7989 2694 8001 2746
rect 8001 2694 8015 2746
rect 8039 2694 8053 2746
rect 8053 2694 8065 2746
rect 8065 2694 8095 2746
rect 8119 2694 8129 2746
rect 8129 2694 8175 2746
rect 7879 2692 7935 2694
rect 7959 2692 8015 2694
rect 8039 2692 8095 2694
rect 8119 2692 8175 2694
rect 6561 2202 6617 2204
rect 6641 2202 6697 2204
rect 6721 2202 6777 2204
rect 6801 2202 6857 2204
rect 6561 2150 6607 2202
rect 6607 2150 6617 2202
rect 6641 2150 6671 2202
rect 6671 2150 6683 2202
rect 6683 2150 6697 2202
rect 6721 2150 6735 2202
rect 6735 2150 6747 2202
rect 6747 2150 6777 2202
rect 6801 2150 6811 2202
rect 6811 2150 6857 2202
rect 6561 2148 6617 2150
rect 6641 2148 6697 2150
rect 6721 2148 6777 2150
rect 6801 2148 6857 2150
rect 8539 2202 8595 2204
rect 8619 2202 8675 2204
rect 8699 2202 8755 2204
rect 8779 2202 8835 2204
rect 8539 2150 8585 2202
rect 8585 2150 8595 2202
rect 8619 2150 8649 2202
rect 8649 2150 8661 2202
rect 8661 2150 8675 2202
rect 8699 2150 8713 2202
rect 8713 2150 8725 2202
rect 8725 2150 8755 2202
rect 8779 2150 8789 2202
rect 8789 2150 8835 2202
rect 8539 2148 8595 2150
rect 8619 2148 8675 2150
rect 8699 2148 8755 2150
rect 8779 2148 8835 2150
<< metal3 >>
rect 2595 9824 2911 9825
rect 2595 9760 2601 9824
rect 2665 9760 2681 9824
rect 2745 9760 2761 9824
rect 2825 9760 2841 9824
rect 2905 9760 2911 9824
rect 2595 9759 2911 9760
rect 4573 9824 4889 9825
rect 4573 9760 4579 9824
rect 4643 9760 4659 9824
rect 4723 9760 4739 9824
rect 4803 9760 4819 9824
rect 4883 9760 4889 9824
rect 4573 9759 4889 9760
rect 6551 9824 6867 9825
rect 6551 9760 6557 9824
rect 6621 9760 6637 9824
rect 6701 9760 6717 9824
rect 6781 9760 6797 9824
rect 6861 9760 6867 9824
rect 6551 9759 6867 9760
rect 8529 9824 8845 9825
rect 8529 9760 8535 9824
rect 8599 9760 8615 9824
rect 8679 9760 8695 9824
rect 8759 9760 8775 9824
rect 8839 9760 8845 9824
rect 8529 9759 8845 9760
rect 1935 9280 2251 9281
rect 1935 9216 1941 9280
rect 2005 9216 2021 9280
rect 2085 9216 2101 9280
rect 2165 9216 2181 9280
rect 2245 9216 2251 9280
rect 1935 9215 2251 9216
rect 3913 9280 4229 9281
rect 3913 9216 3919 9280
rect 3983 9216 3999 9280
rect 4063 9216 4079 9280
rect 4143 9216 4159 9280
rect 4223 9216 4229 9280
rect 3913 9215 4229 9216
rect 5891 9280 6207 9281
rect 5891 9216 5897 9280
rect 5961 9216 5977 9280
rect 6041 9216 6057 9280
rect 6121 9216 6137 9280
rect 6201 9216 6207 9280
rect 5891 9215 6207 9216
rect 7869 9280 8185 9281
rect 7869 9216 7875 9280
rect 7939 9216 7955 9280
rect 8019 9216 8035 9280
rect 8099 9216 8115 9280
rect 8179 9216 8185 9280
rect 7869 9215 8185 9216
rect 0 8938 800 8968
rect 3601 8938 3667 8941
rect 0 8936 3667 8938
rect 0 8880 3606 8936
rect 3662 8880 3667 8936
rect 0 8878 3667 8880
rect 0 8848 800 8878
rect 3601 8875 3667 8878
rect 2595 8736 2911 8737
rect 2595 8672 2601 8736
rect 2665 8672 2681 8736
rect 2745 8672 2761 8736
rect 2825 8672 2841 8736
rect 2905 8672 2911 8736
rect 2595 8671 2911 8672
rect 4573 8736 4889 8737
rect 4573 8672 4579 8736
rect 4643 8672 4659 8736
rect 4723 8672 4739 8736
rect 4803 8672 4819 8736
rect 4883 8672 4889 8736
rect 4573 8671 4889 8672
rect 6551 8736 6867 8737
rect 6551 8672 6557 8736
rect 6621 8672 6637 8736
rect 6701 8672 6717 8736
rect 6781 8672 6797 8736
rect 6861 8672 6867 8736
rect 6551 8671 6867 8672
rect 8529 8736 8845 8737
rect 8529 8672 8535 8736
rect 8599 8672 8615 8736
rect 8679 8672 8695 8736
rect 8759 8672 8775 8736
rect 8839 8672 8845 8736
rect 8529 8671 8845 8672
rect 6361 8394 6427 8397
rect 6318 8392 6427 8394
rect 6318 8336 6366 8392
rect 6422 8336 6427 8392
rect 6318 8331 6427 8336
rect 1935 8192 2251 8193
rect 1935 8128 1941 8192
rect 2005 8128 2021 8192
rect 2085 8128 2101 8192
rect 2165 8128 2181 8192
rect 2245 8128 2251 8192
rect 1935 8127 2251 8128
rect 3913 8192 4229 8193
rect 3913 8128 3919 8192
rect 3983 8128 3999 8192
rect 4063 8128 4079 8192
rect 4143 8128 4159 8192
rect 4223 8128 4229 8192
rect 3913 8127 4229 8128
rect 5891 8192 6207 8193
rect 5891 8128 5897 8192
rect 5961 8128 5977 8192
rect 6041 8128 6057 8192
rect 6121 8128 6137 8192
rect 6201 8128 6207 8192
rect 5891 8127 6207 8128
rect 5901 7986 5967 7989
rect 6318 7986 6378 8331
rect 7869 8192 8185 8193
rect 7869 8128 7875 8192
rect 7939 8128 7955 8192
rect 8019 8128 8035 8192
rect 8099 8128 8115 8192
rect 8179 8128 8185 8192
rect 7869 8127 8185 8128
rect 5901 7984 6378 7986
rect 5901 7928 5906 7984
rect 5962 7928 6378 7984
rect 5901 7926 6378 7928
rect 7557 7986 7623 7989
rect 8109 7986 8175 7989
rect 7557 7984 8175 7986
rect 7557 7928 7562 7984
rect 7618 7928 8114 7984
rect 8170 7928 8175 7984
rect 7557 7926 8175 7928
rect 5901 7923 5967 7926
rect 7557 7923 7623 7926
rect 8109 7923 8175 7926
rect 5073 7850 5139 7853
rect 6361 7850 6427 7853
rect 5073 7848 6427 7850
rect 5073 7792 5078 7848
rect 5134 7792 6366 7848
rect 6422 7792 6427 7848
rect 5073 7790 6427 7792
rect 5073 7787 5139 7790
rect 6361 7787 6427 7790
rect 2595 7648 2911 7649
rect 2595 7584 2601 7648
rect 2665 7584 2681 7648
rect 2745 7584 2761 7648
rect 2825 7584 2841 7648
rect 2905 7584 2911 7648
rect 2595 7583 2911 7584
rect 4573 7648 4889 7649
rect 4573 7584 4579 7648
rect 4643 7584 4659 7648
rect 4723 7584 4739 7648
rect 4803 7584 4819 7648
rect 4883 7584 4889 7648
rect 4573 7583 4889 7584
rect 6551 7648 6867 7649
rect 6551 7584 6557 7648
rect 6621 7584 6637 7648
rect 6701 7584 6717 7648
rect 6781 7584 6797 7648
rect 6861 7584 6867 7648
rect 6551 7583 6867 7584
rect 8529 7648 8845 7649
rect 8529 7584 8535 7648
rect 8599 7584 8615 7648
rect 8679 7584 8695 7648
rect 8759 7584 8775 7648
rect 8839 7584 8845 7648
rect 8529 7583 8845 7584
rect 9029 7578 9095 7581
rect 9412 7578 10212 7608
rect 9029 7576 10212 7578
rect 9029 7520 9034 7576
rect 9090 7520 10212 7576
rect 9029 7518 10212 7520
rect 9029 7515 9095 7518
rect 9412 7488 10212 7518
rect 5625 7306 5691 7309
rect 6085 7306 6151 7309
rect 5625 7304 6151 7306
rect 5625 7248 5630 7304
rect 5686 7248 6090 7304
rect 6146 7248 6151 7304
rect 5625 7246 6151 7248
rect 5625 7243 5691 7246
rect 6085 7243 6151 7246
rect 1935 7104 2251 7105
rect 1935 7040 1941 7104
rect 2005 7040 2021 7104
rect 2085 7040 2101 7104
rect 2165 7040 2181 7104
rect 2245 7040 2251 7104
rect 1935 7039 2251 7040
rect 3913 7104 4229 7105
rect 3913 7040 3919 7104
rect 3983 7040 3999 7104
rect 4063 7040 4079 7104
rect 4143 7040 4159 7104
rect 4223 7040 4229 7104
rect 3913 7039 4229 7040
rect 5891 7104 6207 7105
rect 5891 7040 5897 7104
rect 5961 7040 5977 7104
rect 6041 7040 6057 7104
rect 6121 7040 6137 7104
rect 6201 7040 6207 7104
rect 5891 7039 6207 7040
rect 7869 7104 8185 7105
rect 7869 7040 7875 7104
rect 7939 7040 7955 7104
rect 8019 7040 8035 7104
rect 8099 7040 8115 7104
rect 8179 7040 8185 7104
rect 7869 7039 8185 7040
rect 2595 6560 2911 6561
rect 2595 6496 2601 6560
rect 2665 6496 2681 6560
rect 2745 6496 2761 6560
rect 2825 6496 2841 6560
rect 2905 6496 2911 6560
rect 2595 6495 2911 6496
rect 4573 6560 4889 6561
rect 4573 6496 4579 6560
rect 4643 6496 4659 6560
rect 4723 6496 4739 6560
rect 4803 6496 4819 6560
rect 4883 6496 4889 6560
rect 4573 6495 4889 6496
rect 6551 6560 6867 6561
rect 6551 6496 6557 6560
rect 6621 6496 6637 6560
rect 6701 6496 6717 6560
rect 6781 6496 6797 6560
rect 6861 6496 6867 6560
rect 6551 6495 6867 6496
rect 8529 6560 8845 6561
rect 8529 6496 8535 6560
rect 8599 6496 8615 6560
rect 8679 6496 8695 6560
rect 8759 6496 8775 6560
rect 8839 6496 8845 6560
rect 8529 6495 8845 6496
rect 1761 6354 1827 6357
rect 4521 6354 4587 6357
rect 1761 6352 4587 6354
rect 1761 6296 1766 6352
rect 1822 6296 4526 6352
rect 4582 6296 4587 6352
rect 1761 6294 4587 6296
rect 1761 6291 1827 6294
rect 4521 6291 4587 6294
rect 2865 6218 2931 6221
rect 3877 6218 3943 6221
rect 2865 6216 3943 6218
rect 2865 6160 2870 6216
rect 2926 6160 3882 6216
rect 3938 6160 3943 6216
rect 2865 6158 3943 6160
rect 2865 6155 2931 6158
rect 3877 6155 3943 6158
rect 1935 6016 2251 6017
rect 1935 5952 1941 6016
rect 2005 5952 2021 6016
rect 2085 5952 2101 6016
rect 2165 5952 2181 6016
rect 2245 5952 2251 6016
rect 1935 5951 2251 5952
rect 3913 6016 4229 6017
rect 3913 5952 3919 6016
rect 3983 5952 3999 6016
rect 4063 5952 4079 6016
rect 4143 5952 4159 6016
rect 4223 5952 4229 6016
rect 3913 5951 4229 5952
rect 5891 6016 6207 6017
rect 5891 5952 5897 6016
rect 5961 5952 5977 6016
rect 6041 5952 6057 6016
rect 6121 5952 6137 6016
rect 6201 5952 6207 6016
rect 5891 5951 6207 5952
rect 7869 6016 8185 6017
rect 7869 5952 7875 6016
rect 7939 5952 7955 6016
rect 8019 5952 8035 6016
rect 8099 5952 8115 6016
rect 8179 5952 8185 6016
rect 7869 5951 8185 5952
rect 5165 5946 5231 5949
rect 4478 5944 5231 5946
rect 4478 5888 5170 5944
rect 5226 5888 5231 5944
rect 4478 5886 5231 5888
rect 3877 5810 3943 5813
rect 4478 5810 4538 5886
rect 5165 5883 5231 5886
rect 3877 5808 4538 5810
rect 3877 5752 3882 5808
rect 3938 5752 4538 5808
rect 3877 5750 4538 5752
rect 3877 5747 3943 5750
rect 4153 5674 4219 5677
rect 5533 5674 5599 5677
rect 4153 5672 5599 5674
rect 4153 5616 4158 5672
rect 4214 5616 5538 5672
rect 5594 5616 5599 5672
rect 4153 5614 5599 5616
rect 4153 5611 4219 5614
rect 5533 5611 5599 5614
rect 2595 5472 2911 5473
rect 2595 5408 2601 5472
rect 2665 5408 2681 5472
rect 2745 5408 2761 5472
rect 2825 5408 2841 5472
rect 2905 5408 2911 5472
rect 2595 5407 2911 5408
rect 4573 5472 4889 5473
rect 4573 5408 4579 5472
rect 4643 5408 4659 5472
rect 4723 5408 4739 5472
rect 4803 5408 4819 5472
rect 4883 5408 4889 5472
rect 4573 5407 4889 5408
rect 6551 5472 6867 5473
rect 6551 5408 6557 5472
rect 6621 5408 6637 5472
rect 6701 5408 6717 5472
rect 6781 5408 6797 5472
rect 6861 5408 6867 5472
rect 6551 5407 6867 5408
rect 8529 5472 8845 5473
rect 8529 5408 8535 5472
rect 8599 5408 8615 5472
rect 8679 5408 8695 5472
rect 8759 5408 8775 5472
rect 8839 5408 8845 5472
rect 8529 5407 8845 5408
rect 4981 5402 5047 5405
rect 4981 5400 6378 5402
rect 4981 5344 4986 5400
rect 5042 5344 6378 5400
rect 4981 5342 6378 5344
rect 4981 5339 5047 5342
rect 6318 5266 6378 5342
rect 6453 5266 6519 5269
rect 6318 5264 6519 5266
rect 6318 5208 6458 5264
rect 6514 5208 6519 5264
rect 6318 5206 6519 5208
rect 6453 5203 6519 5206
rect 5165 5130 5231 5133
rect 6085 5130 6151 5133
rect 6637 5130 6703 5133
rect 5165 5128 6703 5130
rect 5165 5072 5170 5128
rect 5226 5072 6090 5128
rect 6146 5072 6642 5128
rect 6698 5072 6703 5128
rect 5165 5070 6703 5072
rect 5165 5067 5231 5070
rect 6085 5067 6151 5070
rect 6637 5067 6703 5070
rect 5073 4994 5139 4997
rect 5625 4994 5691 4997
rect 5073 4992 5691 4994
rect 5073 4936 5078 4992
rect 5134 4936 5630 4992
rect 5686 4936 5691 4992
rect 5073 4934 5691 4936
rect 5073 4931 5139 4934
rect 5625 4931 5691 4934
rect 1935 4928 2251 4929
rect 1935 4864 1941 4928
rect 2005 4864 2021 4928
rect 2085 4864 2101 4928
rect 2165 4864 2181 4928
rect 2245 4864 2251 4928
rect 1935 4863 2251 4864
rect 3913 4928 4229 4929
rect 3913 4864 3919 4928
rect 3983 4864 3999 4928
rect 4063 4864 4079 4928
rect 4143 4864 4159 4928
rect 4223 4864 4229 4928
rect 3913 4863 4229 4864
rect 5891 4928 6207 4929
rect 5891 4864 5897 4928
rect 5961 4864 5977 4928
rect 6041 4864 6057 4928
rect 6121 4864 6137 4928
rect 6201 4864 6207 4928
rect 5891 4863 6207 4864
rect 7869 4928 8185 4929
rect 7869 4864 7875 4928
rect 7939 4864 7955 4928
rect 8019 4864 8035 4928
rect 8099 4864 8115 4928
rect 8179 4864 8185 4928
rect 7869 4863 8185 4864
rect 2865 4858 2931 4861
rect 2454 4856 2931 4858
rect 2454 4800 2870 4856
rect 2926 4800 2931 4856
rect 2454 4798 2931 4800
rect 2129 4722 2195 4725
rect 2454 4722 2514 4798
rect 2865 4795 2931 4798
rect 4613 4858 4679 4861
rect 5257 4858 5323 4861
rect 4613 4856 5323 4858
rect 4613 4800 4618 4856
rect 4674 4800 5262 4856
rect 5318 4800 5323 4856
rect 4613 4798 5323 4800
rect 4613 4795 4679 4798
rect 5257 4795 5323 4798
rect 2129 4720 2514 4722
rect 2129 4664 2134 4720
rect 2190 4664 2514 4720
rect 2129 4662 2514 4664
rect 4797 4722 4863 4725
rect 6453 4722 6519 4725
rect 4797 4720 6519 4722
rect 4797 4664 4802 4720
rect 4858 4664 6458 4720
rect 6514 4664 6519 4720
rect 4797 4662 6519 4664
rect 2129 4659 2195 4662
rect 4797 4659 4863 4662
rect 6453 4659 6519 4662
rect 4061 4586 4127 4589
rect 5993 4586 6059 4589
rect 8569 4586 8635 4589
rect 4061 4584 6059 4586
rect 4061 4528 4066 4584
rect 4122 4528 5998 4584
rect 6054 4528 6059 4584
rect 4061 4526 6059 4528
rect 4061 4523 4127 4526
rect 5993 4523 6059 4526
rect 6134 4584 8635 4586
rect 6134 4528 8574 4584
rect 8630 4528 8635 4584
rect 6134 4526 8635 4528
rect 5257 4450 5323 4453
rect 6134 4450 6194 4526
rect 8569 4523 8635 4526
rect 5257 4448 6194 4450
rect 5257 4392 5262 4448
rect 5318 4392 6194 4448
rect 5257 4390 6194 4392
rect 5257 4387 5323 4390
rect 2595 4384 2911 4385
rect 2595 4320 2601 4384
rect 2665 4320 2681 4384
rect 2745 4320 2761 4384
rect 2825 4320 2841 4384
rect 2905 4320 2911 4384
rect 2595 4319 2911 4320
rect 4573 4384 4889 4385
rect 4573 4320 4579 4384
rect 4643 4320 4659 4384
rect 4723 4320 4739 4384
rect 4803 4320 4819 4384
rect 4883 4320 4889 4384
rect 4573 4319 4889 4320
rect 6551 4384 6867 4385
rect 6551 4320 6557 4384
rect 6621 4320 6637 4384
rect 6701 4320 6717 4384
rect 6781 4320 6797 4384
rect 6861 4320 6867 4384
rect 6551 4319 6867 4320
rect 8529 4384 8845 4385
rect 8529 4320 8535 4384
rect 8599 4320 8615 4384
rect 8679 4320 8695 4384
rect 8759 4320 8775 4384
rect 8839 4320 8845 4384
rect 8529 4319 8845 4320
rect 7005 4314 7071 4317
rect 7005 4312 7114 4314
rect 7005 4256 7010 4312
rect 7066 4256 7114 4312
rect 7005 4251 7114 4256
rect 1761 4042 1827 4045
rect 7054 4042 7114 4251
rect 1761 4040 7114 4042
rect 1761 3984 1766 4040
rect 1822 3984 7114 4040
rect 1761 3982 7114 3984
rect 1761 3979 1827 3982
rect 1935 3840 2251 3841
rect 1935 3776 1941 3840
rect 2005 3776 2021 3840
rect 2085 3776 2101 3840
rect 2165 3776 2181 3840
rect 2245 3776 2251 3840
rect 1935 3775 2251 3776
rect 3913 3840 4229 3841
rect 3913 3776 3919 3840
rect 3983 3776 3999 3840
rect 4063 3776 4079 3840
rect 4143 3776 4159 3840
rect 4223 3776 4229 3840
rect 3913 3775 4229 3776
rect 5891 3840 6207 3841
rect 5891 3776 5897 3840
rect 5961 3776 5977 3840
rect 6041 3776 6057 3840
rect 6121 3776 6137 3840
rect 6201 3776 6207 3840
rect 5891 3775 6207 3776
rect 7869 3840 8185 3841
rect 7869 3776 7875 3840
rect 7939 3776 7955 3840
rect 8019 3776 8035 3840
rect 8099 3776 8115 3840
rect 8179 3776 8185 3840
rect 7869 3775 8185 3776
rect 3969 3634 4035 3637
rect 5165 3634 5231 3637
rect 3969 3632 5231 3634
rect 3969 3576 3974 3632
rect 4030 3576 5170 3632
rect 5226 3576 5231 3632
rect 3969 3574 5231 3576
rect 3969 3571 4035 3574
rect 5165 3571 5231 3574
rect 1485 3498 1551 3501
rect 8017 3498 8083 3501
rect 1485 3496 8083 3498
rect 1485 3440 1490 3496
rect 1546 3440 8022 3496
rect 8078 3440 8083 3496
rect 1485 3438 8083 3440
rect 1485 3435 1551 3438
rect 8017 3435 8083 3438
rect 2595 3296 2911 3297
rect 2595 3232 2601 3296
rect 2665 3232 2681 3296
rect 2745 3232 2761 3296
rect 2825 3232 2841 3296
rect 2905 3232 2911 3296
rect 2595 3231 2911 3232
rect 4573 3296 4889 3297
rect 4573 3232 4579 3296
rect 4643 3232 4659 3296
rect 4723 3232 4739 3296
rect 4803 3232 4819 3296
rect 4883 3232 4889 3296
rect 4573 3231 4889 3232
rect 6551 3296 6867 3297
rect 6551 3232 6557 3296
rect 6621 3232 6637 3296
rect 6701 3232 6717 3296
rect 6781 3232 6797 3296
rect 6861 3232 6867 3296
rect 6551 3231 6867 3232
rect 8529 3296 8845 3297
rect 8529 3232 8535 3296
rect 8599 3232 8615 3296
rect 8679 3232 8695 3296
rect 8759 3232 8775 3296
rect 8839 3232 8845 3296
rect 8529 3231 8845 3232
rect 3233 3090 3299 3093
rect 6913 3090 6979 3093
rect 3233 3088 6979 3090
rect 3233 3032 3238 3088
rect 3294 3032 6918 3088
rect 6974 3032 6979 3088
rect 3233 3030 6979 3032
rect 3233 3027 3299 3030
rect 6913 3027 6979 3030
rect 2037 2954 2103 2957
rect 8385 2954 8451 2957
rect 2037 2952 8451 2954
rect 2037 2896 2042 2952
rect 2098 2896 8390 2952
rect 8446 2896 8451 2952
rect 2037 2894 8451 2896
rect 2037 2891 2103 2894
rect 8385 2891 8451 2894
rect 1935 2752 2251 2753
rect 1935 2688 1941 2752
rect 2005 2688 2021 2752
rect 2085 2688 2101 2752
rect 2165 2688 2181 2752
rect 2245 2688 2251 2752
rect 1935 2687 2251 2688
rect 3913 2752 4229 2753
rect 3913 2688 3919 2752
rect 3983 2688 3999 2752
rect 4063 2688 4079 2752
rect 4143 2688 4159 2752
rect 4223 2688 4229 2752
rect 3913 2687 4229 2688
rect 5891 2752 6207 2753
rect 5891 2688 5897 2752
rect 5961 2688 5977 2752
rect 6041 2688 6057 2752
rect 6121 2688 6137 2752
rect 6201 2688 6207 2752
rect 5891 2687 6207 2688
rect 7869 2752 8185 2753
rect 7869 2688 7875 2752
rect 7939 2688 7955 2752
rect 8019 2688 8035 2752
rect 8099 2688 8115 2752
rect 8179 2688 8185 2752
rect 7869 2687 8185 2688
rect 2497 2546 2563 2549
rect 5073 2546 5139 2549
rect 2497 2544 5139 2546
rect 2497 2488 2502 2544
rect 2558 2488 5078 2544
rect 5134 2488 5139 2544
rect 2497 2486 5139 2488
rect 2497 2483 2563 2486
rect 5073 2483 5139 2486
rect 3417 2410 3483 2413
rect 5625 2410 5691 2413
rect 3417 2408 5691 2410
rect 3417 2352 3422 2408
rect 3478 2352 5630 2408
rect 5686 2352 5691 2408
rect 3417 2350 5691 2352
rect 3417 2347 3483 2350
rect 5625 2347 5691 2350
rect 2595 2208 2911 2209
rect 2595 2144 2601 2208
rect 2665 2144 2681 2208
rect 2745 2144 2761 2208
rect 2825 2144 2841 2208
rect 2905 2144 2911 2208
rect 2595 2143 2911 2144
rect 4573 2208 4889 2209
rect 4573 2144 4579 2208
rect 4643 2144 4659 2208
rect 4723 2144 4739 2208
rect 4803 2144 4819 2208
rect 4883 2144 4889 2208
rect 4573 2143 4889 2144
rect 6551 2208 6867 2209
rect 6551 2144 6557 2208
rect 6621 2144 6637 2208
rect 6701 2144 6717 2208
rect 6781 2144 6797 2208
rect 6861 2144 6867 2208
rect 6551 2143 6867 2144
rect 8529 2208 8845 2209
rect 8529 2144 8535 2208
rect 8599 2144 8615 2208
rect 8679 2144 8695 2208
rect 8759 2144 8775 2208
rect 8839 2144 8845 2208
rect 8529 2143 8845 2144
<< via3 >>
rect 2601 9820 2665 9824
rect 2601 9764 2605 9820
rect 2605 9764 2661 9820
rect 2661 9764 2665 9820
rect 2601 9760 2665 9764
rect 2681 9820 2745 9824
rect 2681 9764 2685 9820
rect 2685 9764 2741 9820
rect 2741 9764 2745 9820
rect 2681 9760 2745 9764
rect 2761 9820 2825 9824
rect 2761 9764 2765 9820
rect 2765 9764 2821 9820
rect 2821 9764 2825 9820
rect 2761 9760 2825 9764
rect 2841 9820 2905 9824
rect 2841 9764 2845 9820
rect 2845 9764 2901 9820
rect 2901 9764 2905 9820
rect 2841 9760 2905 9764
rect 4579 9820 4643 9824
rect 4579 9764 4583 9820
rect 4583 9764 4639 9820
rect 4639 9764 4643 9820
rect 4579 9760 4643 9764
rect 4659 9820 4723 9824
rect 4659 9764 4663 9820
rect 4663 9764 4719 9820
rect 4719 9764 4723 9820
rect 4659 9760 4723 9764
rect 4739 9820 4803 9824
rect 4739 9764 4743 9820
rect 4743 9764 4799 9820
rect 4799 9764 4803 9820
rect 4739 9760 4803 9764
rect 4819 9820 4883 9824
rect 4819 9764 4823 9820
rect 4823 9764 4879 9820
rect 4879 9764 4883 9820
rect 4819 9760 4883 9764
rect 6557 9820 6621 9824
rect 6557 9764 6561 9820
rect 6561 9764 6617 9820
rect 6617 9764 6621 9820
rect 6557 9760 6621 9764
rect 6637 9820 6701 9824
rect 6637 9764 6641 9820
rect 6641 9764 6697 9820
rect 6697 9764 6701 9820
rect 6637 9760 6701 9764
rect 6717 9820 6781 9824
rect 6717 9764 6721 9820
rect 6721 9764 6777 9820
rect 6777 9764 6781 9820
rect 6717 9760 6781 9764
rect 6797 9820 6861 9824
rect 6797 9764 6801 9820
rect 6801 9764 6857 9820
rect 6857 9764 6861 9820
rect 6797 9760 6861 9764
rect 8535 9820 8599 9824
rect 8535 9764 8539 9820
rect 8539 9764 8595 9820
rect 8595 9764 8599 9820
rect 8535 9760 8599 9764
rect 8615 9820 8679 9824
rect 8615 9764 8619 9820
rect 8619 9764 8675 9820
rect 8675 9764 8679 9820
rect 8615 9760 8679 9764
rect 8695 9820 8759 9824
rect 8695 9764 8699 9820
rect 8699 9764 8755 9820
rect 8755 9764 8759 9820
rect 8695 9760 8759 9764
rect 8775 9820 8839 9824
rect 8775 9764 8779 9820
rect 8779 9764 8835 9820
rect 8835 9764 8839 9820
rect 8775 9760 8839 9764
rect 1941 9276 2005 9280
rect 1941 9220 1945 9276
rect 1945 9220 2001 9276
rect 2001 9220 2005 9276
rect 1941 9216 2005 9220
rect 2021 9276 2085 9280
rect 2021 9220 2025 9276
rect 2025 9220 2081 9276
rect 2081 9220 2085 9276
rect 2021 9216 2085 9220
rect 2101 9276 2165 9280
rect 2101 9220 2105 9276
rect 2105 9220 2161 9276
rect 2161 9220 2165 9276
rect 2101 9216 2165 9220
rect 2181 9276 2245 9280
rect 2181 9220 2185 9276
rect 2185 9220 2241 9276
rect 2241 9220 2245 9276
rect 2181 9216 2245 9220
rect 3919 9276 3983 9280
rect 3919 9220 3923 9276
rect 3923 9220 3979 9276
rect 3979 9220 3983 9276
rect 3919 9216 3983 9220
rect 3999 9276 4063 9280
rect 3999 9220 4003 9276
rect 4003 9220 4059 9276
rect 4059 9220 4063 9276
rect 3999 9216 4063 9220
rect 4079 9276 4143 9280
rect 4079 9220 4083 9276
rect 4083 9220 4139 9276
rect 4139 9220 4143 9276
rect 4079 9216 4143 9220
rect 4159 9276 4223 9280
rect 4159 9220 4163 9276
rect 4163 9220 4219 9276
rect 4219 9220 4223 9276
rect 4159 9216 4223 9220
rect 5897 9276 5961 9280
rect 5897 9220 5901 9276
rect 5901 9220 5957 9276
rect 5957 9220 5961 9276
rect 5897 9216 5961 9220
rect 5977 9276 6041 9280
rect 5977 9220 5981 9276
rect 5981 9220 6037 9276
rect 6037 9220 6041 9276
rect 5977 9216 6041 9220
rect 6057 9276 6121 9280
rect 6057 9220 6061 9276
rect 6061 9220 6117 9276
rect 6117 9220 6121 9276
rect 6057 9216 6121 9220
rect 6137 9276 6201 9280
rect 6137 9220 6141 9276
rect 6141 9220 6197 9276
rect 6197 9220 6201 9276
rect 6137 9216 6201 9220
rect 7875 9276 7939 9280
rect 7875 9220 7879 9276
rect 7879 9220 7935 9276
rect 7935 9220 7939 9276
rect 7875 9216 7939 9220
rect 7955 9276 8019 9280
rect 7955 9220 7959 9276
rect 7959 9220 8015 9276
rect 8015 9220 8019 9276
rect 7955 9216 8019 9220
rect 8035 9276 8099 9280
rect 8035 9220 8039 9276
rect 8039 9220 8095 9276
rect 8095 9220 8099 9276
rect 8035 9216 8099 9220
rect 8115 9276 8179 9280
rect 8115 9220 8119 9276
rect 8119 9220 8175 9276
rect 8175 9220 8179 9276
rect 8115 9216 8179 9220
rect 2601 8732 2665 8736
rect 2601 8676 2605 8732
rect 2605 8676 2661 8732
rect 2661 8676 2665 8732
rect 2601 8672 2665 8676
rect 2681 8732 2745 8736
rect 2681 8676 2685 8732
rect 2685 8676 2741 8732
rect 2741 8676 2745 8732
rect 2681 8672 2745 8676
rect 2761 8732 2825 8736
rect 2761 8676 2765 8732
rect 2765 8676 2821 8732
rect 2821 8676 2825 8732
rect 2761 8672 2825 8676
rect 2841 8732 2905 8736
rect 2841 8676 2845 8732
rect 2845 8676 2901 8732
rect 2901 8676 2905 8732
rect 2841 8672 2905 8676
rect 4579 8732 4643 8736
rect 4579 8676 4583 8732
rect 4583 8676 4639 8732
rect 4639 8676 4643 8732
rect 4579 8672 4643 8676
rect 4659 8732 4723 8736
rect 4659 8676 4663 8732
rect 4663 8676 4719 8732
rect 4719 8676 4723 8732
rect 4659 8672 4723 8676
rect 4739 8732 4803 8736
rect 4739 8676 4743 8732
rect 4743 8676 4799 8732
rect 4799 8676 4803 8732
rect 4739 8672 4803 8676
rect 4819 8732 4883 8736
rect 4819 8676 4823 8732
rect 4823 8676 4879 8732
rect 4879 8676 4883 8732
rect 4819 8672 4883 8676
rect 6557 8732 6621 8736
rect 6557 8676 6561 8732
rect 6561 8676 6617 8732
rect 6617 8676 6621 8732
rect 6557 8672 6621 8676
rect 6637 8732 6701 8736
rect 6637 8676 6641 8732
rect 6641 8676 6697 8732
rect 6697 8676 6701 8732
rect 6637 8672 6701 8676
rect 6717 8732 6781 8736
rect 6717 8676 6721 8732
rect 6721 8676 6777 8732
rect 6777 8676 6781 8732
rect 6717 8672 6781 8676
rect 6797 8732 6861 8736
rect 6797 8676 6801 8732
rect 6801 8676 6857 8732
rect 6857 8676 6861 8732
rect 6797 8672 6861 8676
rect 8535 8732 8599 8736
rect 8535 8676 8539 8732
rect 8539 8676 8595 8732
rect 8595 8676 8599 8732
rect 8535 8672 8599 8676
rect 8615 8732 8679 8736
rect 8615 8676 8619 8732
rect 8619 8676 8675 8732
rect 8675 8676 8679 8732
rect 8615 8672 8679 8676
rect 8695 8732 8759 8736
rect 8695 8676 8699 8732
rect 8699 8676 8755 8732
rect 8755 8676 8759 8732
rect 8695 8672 8759 8676
rect 8775 8732 8839 8736
rect 8775 8676 8779 8732
rect 8779 8676 8835 8732
rect 8835 8676 8839 8732
rect 8775 8672 8839 8676
rect 1941 8188 2005 8192
rect 1941 8132 1945 8188
rect 1945 8132 2001 8188
rect 2001 8132 2005 8188
rect 1941 8128 2005 8132
rect 2021 8188 2085 8192
rect 2021 8132 2025 8188
rect 2025 8132 2081 8188
rect 2081 8132 2085 8188
rect 2021 8128 2085 8132
rect 2101 8188 2165 8192
rect 2101 8132 2105 8188
rect 2105 8132 2161 8188
rect 2161 8132 2165 8188
rect 2101 8128 2165 8132
rect 2181 8188 2245 8192
rect 2181 8132 2185 8188
rect 2185 8132 2241 8188
rect 2241 8132 2245 8188
rect 2181 8128 2245 8132
rect 3919 8188 3983 8192
rect 3919 8132 3923 8188
rect 3923 8132 3979 8188
rect 3979 8132 3983 8188
rect 3919 8128 3983 8132
rect 3999 8188 4063 8192
rect 3999 8132 4003 8188
rect 4003 8132 4059 8188
rect 4059 8132 4063 8188
rect 3999 8128 4063 8132
rect 4079 8188 4143 8192
rect 4079 8132 4083 8188
rect 4083 8132 4139 8188
rect 4139 8132 4143 8188
rect 4079 8128 4143 8132
rect 4159 8188 4223 8192
rect 4159 8132 4163 8188
rect 4163 8132 4219 8188
rect 4219 8132 4223 8188
rect 4159 8128 4223 8132
rect 5897 8188 5961 8192
rect 5897 8132 5901 8188
rect 5901 8132 5957 8188
rect 5957 8132 5961 8188
rect 5897 8128 5961 8132
rect 5977 8188 6041 8192
rect 5977 8132 5981 8188
rect 5981 8132 6037 8188
rect 6037 8132 6041 8188
rect 5977 8128 6041 8132
rect 6057 8188 6121 8192
rect 6057 8132 6061 8188
rect 6061 8132 6117 8188
rect 6117 8132 6121 8188
rect 6057 8128 6121 8132
rect 6137 8188 6201 8192
rect 6137 8132 6141 8188
rect 6141 8132 6197 8188
rect 6197 8132 6201 8188
rect 6137 8128 6201 8132
rect 7875 8188 7939 8192
rect 7875 8132 7879 8188
rect 7879 8132 7935 8188
rect 7935 8132 7939 8188
rect 7875 8128 7939 8132
rect 7955 8188 8019 8192
rect 7955 8132 7959 8188
rect 7959 8132 8015 8188
rect 8015 8132 8019 8188
rect 7955 8128 8019 8132
rect 8035 8188 8099 8192
rect 8035 8132 8039 8188
rect 8039 8132 8095 8188
rect 8095 8132 8099 8188
rect 8035 8128 8099 8132
rect 8115 8188 8179 8192
rect 8115 8132 8119 8188
rect 8119 8132 8175 8188
rect 8175 8132 8179 8188
rect 8115 8128 8179 8132
rect 2601 7644 2665 7648
rect 2601 7588 2605 7644
rect 2605 7588 2661 7644
rect 2661 7588 2665 7644
rect 2601 7584 2665 7588
rect 2681 7644 2745 7648
rect 2681 7588 2685 7644
rect 2685 7588 2741 7644
rect 2741 7588 2745 7644
rect 2681 7584 2745 7588
rect 2761 7644 2825 7648
rect 2761 7588 2765 7644
rect 2765 7588 2821 7644
rect 2821 7588 2825 7644
rect 2761 7584 2825 7588
rect 2841 7644 2905 7648
rect 2841 7588 2845 7644
rect 2845 7588 2901 7644
rect 2901 7588 2905 7644
rect 2841 7584 2905 7588
rect 4579 7644 4643 7648
rect 4579 7588 4583 7644
rect 4583 7588 4639 7644
rect 4639 7588 4643 7644
rect 4579 7584 4643 7588
rect 4659 7644 4723 7648
rect 4659 7588 4663 7644
rect 4663 7588 4719 7644
rect 4719 7588 4723 7644
rect 4659 7584 4723 7588
rect 4739 7644 4803 7648
rect 4739 7588 4743 7644
rect 4743 7588 4799 7644
rect 4799 7588 4803 7644
rect 4739 7584 4803 7588
rect 4819 7644 4883 7648
rect 4819 7588 4823 7644
rect 4823 7588 4879 7644
rect 4879 7588 4883 7644
rect 4819 7584 4883 7588
rect 6557 7644 6621 7648
rect 6557 7588 6561 7644
rect 6561 7588 6617 7644
rect 6617 7588 6621 7644
rect 6557 7584 6621 7588
rect 6637 7644 6701 7648
rect 6637 7588 6641 7644
rect 6641 7588 6697 7644
rect 6697 7588 6701 7644
rect 6637 7584 6701 7588
rect 6717 7644 6781 7648
rect 6717 7588 6721 7644
rect 6721 7588 6777 7644
rect 6777 7588 6781 7644
rect 6717 7584 6781 7588
rect 6797 7644 6861 7648
rect 6797 7588 6801 7644
rect 6801 7588 6857 7644
rect 6857 7588 6861 7644
rect 6797 7584 6861 7588
rect 8535 7644 8599 7648
rect 8535 7588 8539 7644
rect 8539 7588 8595 7644
rect 8595 7588 8599 7644
rect 8535 7584 8599 7588
rect 8615 7644 8679 7648
rect 8615 7588 8619 7644
rect 8619 7588 8675 7644
rect 8675 7588 8679 7644
rect 8615 7584 8679 7588
rect 8695 7644 8759 7648
rect 8695 7588 8699 7644
rect 8699 7588 8755 7644
rect 8755 7588 8759 7644
rect 8695 7584 8759 7588
rect 8775 7644 8839 7648
rect 8775 7588 8779 7644
rect 8779 7588 8835 7644
rect 8835 7588 8839 7644
rect 8775 7584 8839 7588
rect 1941 7100 2005 7104
rect 1941 7044 1945 7100
rect 1945 7044 2001 7100
rect 2001 7044 2005 7100
rect 1941 7040 2005 7044
rect 2021 7100 2085 7104
rect 2021 7044 2025 7100
rect 2025 7044 2081 7100
rect 2081 7044 2085 7100
rect 2021 7040 2085 7044
rect 2101 7100 2165 7104
rect 2101 7044 2105 7100
rect 2105 7044 2161 7100
rect 2161 7044 2165 7100
rect 2101 7040 2165 7044
rect 2181 7100 2245 7104
rect 2181 7044 2185 7100
rect 2185 7044 2241 7100
rect 2241 7044 2245 7100
rect 2181 7040 2245 7044
rect 3919 7100 3983 7104
rect 3919 7044 3923 7100
rect 3923 7044 3979 7100
rect 3979 7044 3983 7100
rect 3919 7040 3983 7044
rect 3999 7100 4063 7104
rect 3999 7044 4003 7100
rect 4003 7044 4059 7100
rect 4059 7044 4063 7100
rect 3999 7040 4063 7044
rect 4079 7100 4143 7104
rect 4079 7044 4083 7100
rect 4083 7044 4139 7100
rect 4139 7044 4143 7100
rect 4079 7040 4143 7044
rect 4159 7100 4223 7104
rect 4159 7044 4163 7100
rect 4163 7044 4219 7100
rect 4219 7044 4223 7100
rect 4159 7040 4223 7044
rect 5897 7100 5961 7104
rect 5897 7044 5901 7100
rect 5901 7044 5957 7100
rect 5957 7044 5961 7100
rect 5897 7040 5961 7044
rect 5977 7100 6041 7104
rect 5977 7044 5981 7100
rect 5981 7044 6037 7100
rect 6037 7044 6041 7100
rect 5977 7040 6041 7044
rect 6057 7100 6121 7104
rect 6057 7044 6061 7100
rect 6061 7044 6117 7100
rect 6117 7044 6121 7100
rect 6057 7040 6121 7044
rect 6137 7100 6201 7104
rect 6137 7044 6141 7100
rect 6141 7044 6197 7100
rect 6197 7044 6201 7100
rect 6137 7040 6201 7044
rect 7875 7100 7939 7104
rect 7875 7044 7879 7100
rect 7879 7044 7935 7100
rect 7935 7044 7939 7100
rect 7875 7040 7939 7044
rect 7955 7100 8019 7104
rect 7955 7044 7959 7100
rect 7959 7044 8015 7100
rect 8015 7044 8019 7100
rect 7955 7040 8019 7044
rect 8035 7100 8099 7104
rect 8035 7044 8039 7100
rect 8039 7044 8095 7100
rect 8095 7044 8099 7100
rect 8035 7040 8099 7044
rect 8115 7100 8179 7104
rect 8115 7044 8119 7100
rect 8119 7044 8175 7100
rect 8175 7044 8179 7100
rect 8115 7040 8179 7044
rect 2601 6556 2665 6560
rect 2601 6500 2605 6556
rect 2605 6500 2661 6556
rect 2661 6500 2665 6556
rect 2601 6496 2665 6500
rect 2681 6556 2745 6560
rect 2681 6500 2685 6556
rect 2685 6500 2741 6556
rect 2741 6500 2745 6556
rect 2681 6496 2745 6500
rect 2761 6556 2825 6560
rect 2761 6500 2765 6556
rect 2765 6500 2821 6556
rect 2821 6500 2825 6556
rect 2761 6496 2825 6500
rect 2841 6556 2905 6560
rect 2841 6500 2845 6556
rect 2845 6500 2901 6556
rect 2901 6500 2905 6556
rect 2841 6496 2905 6500
rect 4579 6556 4643 6560
rect 4579 6500 4583 6556
rect 4583 6500 4639 6556
rect 4639 6500 4643 6556
rect 4579 6496 4643 6500
rect 4659 6556 4723 6560
rect 4659 6500 4663 6556
rect 4663 6500 4719 6556
rect 4719 6500 4723 6556
rect 4659 6496 4723 6500
rect 4739 6556 4803 6560
rect 4739 6500 4743 6556
rect 4743 6500 4799 6556
rect 4799 6500 4803 6556
rect 4739 6496 4803 6500
rect 4819 6556 4883 6560
rect 4819 6500 4823 6556
rect 4823 6500 4879 6556
rect 4879 6500 4883 6556
rect 4819 6496 4883 6500
rect 6557 6556 6621 6560
rect 6557 6500 6561 6556
rect 6561 6500 6617 6556
rect 6617 6500 6621 6556
rect 6557 6496 6621 6500
rect 6637 6556 6701 6560
rect 6637 6500 6641 6556
rect 6641 6500 6697 6556
rect 6697 6500 6701 6556
rect 6637 6496 6701 6500
rect 6717 6556 6781 6560
rect 6717 6500 6721 6556
rect 6721 6500 6777 6556
rect 6777 6500 6781 6556
rect 6717 6496 6781 6500
rect 6797 6556 6861 6560
rect 6797 6500 6801 6556
rect 6801 6500 6857 6556
rect 6857 6500 6861 6556
rect 6797 6496 6861 6500
rect 8535 6556 8599 6560
rect 8535 6500 8539 6556
rect 8539 6500 8595 6556
rect 8595 6500 8599 6556
rect 8535 6496 8599 6500
rect 8615 6556 8679 6560
rect 8615 6500 8619 6556
rect 8619 6500 8675 6556
rect 8675 6500 8679 6556
rect 8615 6496 8679 6500
rect 8695 6556 8759 6560
rect 8695 6500 8699 6556
rect 8699 6500 8755 6556
rect 8755 6500 8759 6556
rect 8695 6496 8759 6500
rect 8775 6556 8839 6560
rect 8775 6500 8779 6556
rect 8779 6500 8835 6556
rect 8835 6500 8839 6556
rect 8775 6496 8839 6500
rect 1941 6012 2005 6016
rect 1941 5956 1945 6012
rect 1945 5956 2001 6012
rect 2001 5956 2005 6012
rect 1941 5952 2005 5956
rect 2021 6012 2085 6016
rect 2021 5956 2025 6012
rect 2025 5956 2081 6012
rect 2081 5956 2085 6012
rect 2021 5952 2085 5956
rect 2101 6012 2165 6016
rect 2101 5956 2105 6012
rect 2105 5956 2161 6012
rect 2161 5956 2165 6012
rect 2101 5952 2165 5956
rect 2181 6012 2245 6016
rect 2181 5956 2185 6012
rect 2185 5956 2241 6012
rect 2241 5956 2245 6012
rect 2181 5952 2245 5956
rect 3919 6012 3983 6016
rect 3919 5956 3923 6012
rect 3923 5956 3979 6012
rect 3979 5956 3983 6012
rect 3919 5952 3983 5956
rect 3999 6012 4063 6016
rect 3999 5956 4003 6012
rect 4003 5956 4059 6012
rect 4059 5956 4063 6012
rect 3999 5952 4063 5956
rect 4079 6012 4143 6016
rect 4079 5956 4083 6012
rect 4083 5956 4139 6012
rect 4139 5956 4143 6012
rect 4079 5952 4143 5956
rect 4159 6012 4223 6016
rect 4159 5956 4163 6012
rect 4163 5956 4219 6012
rect 4219 5956 4223 6012
rect 4159 5952 4223 5956
rect 5897 6012 5961 6016
rect 5897 5956 5901 6012
rect 5901 5956 5957 6012
rect 5957 5956 5961 6012
rect 5897 5952 5961 5956
rect 5977 6012 6041 6016
rect 5977 5956 5981 6012
rect 5981 5956 6037 6012
rect 6037 5956 6041 6012
rect 5977 5952 6041 5956
rect 6057 6012 6121 6016
rect 6057 5956 6061 6012
rect 6061 5956 6117 6012
rect 6117 5956 6121 6012
rect 6057 5952 6121 5956
rect 6137 6012 6201 6016
rect 6137 5956 6141 6012
rect 6141 5956 6197 6012
rect 6197 5956 6201 6012
rect 6137 5952 6201 5956
rect 7875 6012 7939 6016
rect 7875 5956 7879 6012
rect 7879 5956 7935 6012
rect 7935 5956 7939 6012
rect 7875 5952 7939 5956
rect 7955 6012 8019 6016
rect 7955 5956 7959 6012
rect 7959 5956 8015 6012
rect 8015 5956 8019 6012
rect 7955 5952 8019 5956
rect 8035 6012 8099 6016
rect 8035 5956 8039 6012
rect 8039 5956 8095 6012
rect 8095 5956 8099 6012
rect 8035 5952 8099 5956
rect 8115 6012 8179 6016
rect 8115 5956 8119 6012
rect 8119 5956 8175 6012
rect 8175 5956 8179 6012
rect 8115 5952 8179 5956
rect 2601 5468 2665 5472
rect 2601 5412 2605 5468
rect 2605 5412 2661 5468
rect 2661 5412 2665 5468
rect 2601 5408 2665 5412
rect 2681 5468 2745 5472
rect 2681 5412 2685 5468
rect 2685 5412 2741 5468
rect 2741 5412 2745 5468
rect 2681 5408 2745 5412
rect 2761 5468 2825 5472
rect 2761 5412 2765 5468
rect 2765 5412 2821 5468
rect 2821 5412 2825 5468
rect 2761 5408 2825 5412
rect 2841 5468 2905 5472
rect 2841 5412 2845 5468
rect 2845 5412 2901 5468
rect 2901 5412 2905 5468
rect 2841 5408 2905 5412
rect 4579 5468 4643 5472
rect 4579 5412 4583 5468
rect 4583 5412 4639 5468
rect 4639 5412 4643 5468
rect 4579 5408 4643 5412
rect 4659 5468 4723 5472
rect 4659 5412 4663 5468
rect 4663 5412 4719 5468
rect 4719 5412 4723 5468
rect 4659 5408 4723 5412
rect 4739 5468 4803 5472
rect 4739 5412 4743 5468
rect 4743 5412 4799 5468
rect 4799 5412 4803 5468
rect 4739 5408 4803 5412
rect 4819 5468 4883 5472
rect 4819 5412 4823 5468
rect 4823 5412 4879 5468
rect 4879 5412 4883 5468
rect 4819 5408 4883 5412
rect 6557 5468 6621 5472
rect 6557 5412 6561 5468
rect 6561 5412 6617 5468
rect 6617 5412 6621 5468
rect 6557 5408 6621 5412
rect 6637 5468 6701 5472
rect 6637 5412 6641 5468
rect 6641 5412 6697 5468
rect 6697 5412 6701 5468
rect 6637 5408 6701 5412
rect 6717 5468 6781 5472
rect 6717 5412 6721 5468
rect 6721 5412 6777 5468
rect 6777 5412 6781 5468
rect 6717 5408 6781 5412
rect 6797 5468 6861 5472
rect 6797 5412 6801 5468
rect 6801 5412 6857 5468
rect 6857 5412 6861 5468
rect 6797 5408 6861 5412
rect 8535 5468 8599 5472
rect 8535 5412 8539 5468
rect 8539 5412 8595 5468
rect 8595 5412 8599 5468
rect 8535 5408 8599 5412
rect 8615 5468 8679 5472
rect 8615 5412 8619 5468
rect 8619 5412 8675 5468
rect 8675 5412 8679 5468
rect 8615 5408 8679 5412
rect 8695 5468 8759 5472
rect 8695 5412 8699 5468
rect 8699 5412 8755 5468
rect 8755 5412 8759 5468
rect 8695 5408 8759 5412
rect 8775 5468 8839 5472
rect 8775 5412 8779 5468
rect 8779 5412 8835 5468
rect 8835 5412 8839 5468
rect 8775 5408 8839 5412
rect 1941 4924 2005 4928
rect 1941 4868 1945 4924
rect 1945 4868 2001 4924
rect 2001 4868 2005 4924
rect 1941 4864 2005 4868
rect 2021 4924 2085 4928
rect 2021 4868 2025 4924
rect 2025 4868 2081 4924
rect 2081 4868 2085 4924
rect 2021 4864 2085 4868
rect 2101 4924 2165 4928
rect 2101 4868 2105 4924
rect 2105 4868 2161 4924
rect 2161 4868 2165 4924
rect 2101 4864 2165 4868
rect 2181 4924 2245 4928
rect 2181 4868 2185 4924
rect 2185 4868 2241 4924
rect 2241 4868 2245 4924
rect 2181 4864 2245 4868
rect 3919 4924 3983 4928
rect 3919 4868 3923 4924
rect 3923 4868 3979 4924
rect 3979 4868 3983 4924
rect 3919 4864 3983 4868
rect 3999 4924 4063 4928
rect 3999 4868 4003 4924
rect 4003 4868 4059 4924
rect 4059 4868 4063 4924
rect 3999 4864 4063 4868
rect 4079 4924 4143 4928
rect 4079 4868 4083 4924
rect 4083 4868 4139 4924
rect 4139 4868 4143 4924
rect 4079 4864 4143 4868
rect 4159 4924 4223 4928
rect 4159 4868 4163 4924
rect 4163 4868 4219 4924
rect 4219 4868 4223 4924
rect 4159 4864 4223 4868
rect 5897 4924 5961 4928
rect 5897 4868 5901 4924
rect 5901 4868 5957 4924
rect 5957 4868 5961 4924
rect 5897 4864 5961 4868
rect 5977 4924 6041 4928
rect 5977 4868 5981 4924
rect 5981 4868 6037 4924
rect 6037 4868 6041 4924
rect 5977 4864 6041 4868
rect 6057 4924 6121 4928
rect 6057 4868 6061 4924
rect 6061 4868 6117 4924
rect 6117 4868 6121 4924
rect 6057 4864 6121 4868
rect 6137 4924 6201 4928
rect 6137 4868 6141 4924
rect 6141 4868 6197 4924
rect 6197 4868 6201 4924
rect 6137 4864 6201 4868
rect 7875 4924 7939 4928
rect 7875 4868 7879 4924
rect 7879 4868 7935 4924
rect 7935 4868 7939 4924
rect 7875 4864 7939 4868
rect 7955 4924 8019 4928
rect 7955 4868 7959 4924
rect 7959 4868 8015 4924
rect 8015 4868 8019 4924
rect 7955 4864 8019 4868
rect 8035 4924 8099 4928
rect 8035 4868 8039 4924
rect 8039 4868 8095 4924
rect 8095 4868 8099 4924
rect 8035 4864 8099 4868
rect 8115 4924 8179 4928
rect 8115 4868 8119 4924
rect 8119 4868 8175 4924
rect 8175 4868 8179 4924
rect 8115 4864 8179 4868
rect 2601 4380 2665 4384
rect 2601 4324 2605 4380
rect 2605 4324 2661 4380
rect 2661 4324 2665 4380
rect 2601 4320 2665 4324
rect 2681 4380 2745 4384
rect 2681 4324 2685 4380
rect 2685 4324 2741 4380
rect 2741 4324 2745 4380
rect 2681 4320 2745 4324
rect 2761 4380 2825 4384
rect 2761 4324 2765 4380
rect 2765 4324 2821 4380
rect 2821 4324 2825 4380
rect 2761 4320 2825 4324
rect 2841 4380 2905 4384
rect 2841 4324 2845 4380
rect 2845 4324 2901 4380
rect 2901 4324 2905 4380
rect 2841 4320 2905 4324
rect 4579 4380 4643 4384
rect 4579 4324 4583 4380
rect 4583 4324 4639 4380
rect 4639 4324 4643 4380
rect 4579 4320 4643 4324
rect 4659 4380 4723 4384
rect 4659 4324 4663 4380
rect 4663 4324 4719 4380
rect 4719 4324 4723 4380
rect 4659 4320 4723 4324
rect 4739 4380 4803 4384
rect 4739 4324 4743 4380
rect 4743 4324 4799 4380
rect 4799 4324 4803 4380
rect 4739 4320 4803 4324
rect 4819 4380 4883 4384
rect 4819 4324 4823 4380
rect 4823 4324 4879 4380
rect 4879 4324 4883 4380
rect 4819 4320 4883 4324
rect 6557 4380 6621 4384
rect 6557 4324 6561 4380
rect 6561 4324 6617 4380
rect 6617 4324 6621 4380
rect 6557 4320 6621 4324
rect 6637 4380 6701 4384
rect 6637 4324 6641 4380
rect 6641 4324 6697 4380
rect 6697 4324 6701 4380
rect 6637 4320 6701 4324
rect 6717 4380 6781 4384
rect 6717 4324 6721 4380
rect 6721 4324 6777 4380
rect 6777 4324 6781 4380
rect 6717 4320 6781 4324
rect 6797 4380 6861 4384
rect 6797 4324 6801 4380
rect 6801 4324 6857 4380
rect 6857 4324 6861 4380
rect 6797 4320 6861 4324
rect 8535 4380 8599 4384
rect 8535 4324 8539 4380
rect 8539 4324 8595 4380
rect 8595 4324 8599 4380
rect 8535 4320 8599 4324
rect 8615 4380 8679 4384
rect 8615 4324 8619 4380
rect 8619 4324 8675 4380
rect 8675 4324 8679 4380
rect 8615 4320 8679 4324
rect 8695 4380 8759 4384
rect 8695 4324 8699 4380
rect 8699 4324 8755 4380
rect 8755 4324 8759 4380
rect 8695 4320 8759 4324
rect 8775 4380 8839 4384
rect 8775 4324 8779 4380
rect 8779 4324 8835 4380
rect 8835 4324 8839 4380
rect 8775 4320 8839 4324
rect 1941 3836 2005 3840
rect 1941 3780 1945 3836
rect 1945 3780 2001 3836
rect 2001 3780 2005 3836
rect 1941 3776 2005 3780
rect 2021 3836 2085 3840
rect 2021 3780 2025 3836
rect 2025 3780 2081 3836
rect 2081 3780 2085 3836
rect 2021 3776 2085 3780
rect 2101 3836 2165 3840
rect 2101 3780 2105 3836
rect 2105 3780 2161 3836
rect 2161 3780 2165 3836
rect 2101 3776 2165 3780
rect 2181 3836 2245 3840
rect 2181 3780 2185 3836
rect 2185 3780 2241 3836
rect 2241 3780 2245 3836
rect 2181 3776 2245 3780
rect 3919 3836 3983 3840
rect 3919 3780 3923 3836
rect 3923 3780 3979 3836
rect 3979 3780 3983 3836
rect 3919 3776 3983 3780
rect 3999 3836 4063 3840
rect 3999 3780 4003 3836
rect 4003 3780 4059 3836
rect 4059 3780 4063 3836
rect 3999 3776 4063 3780
rect 4079 3836 4143 3840
rect 4079 3780 4083 3836
rect 4083 3780 4139 3836
rect 4139 3780 4143 3836
rect 4079 3776 4143 3780
rect 4159 3836 4223 3840
rect 4159 3780 4163 3836
rect 4163 3780 4219 3836
rect 4219 3780 4223 3836
rect 4159 3776 4223 3780
rect 5897 3836 5961 3840
rect 5897 3780 5901 3836
rect 5901 3780 5957 3836
rect 5957 3780 5961 3836
rect 5897 3776 5961 3780
rect 5977 3836 6041 3840
rect 5977 3780 5981 3836
rect 5981 3780 6037 3836
rect 6037 3780 6041 3836
rect 5977 3776 6041 3780
rect 6057 3836 6121 3840
rect 6057 3780 6061 3836
rect 6061 3780 6117 3836
rect 6117 3780 6121 3836
rect 6057 3776 6121 3780
rect 6137 3836 6201 3840
rect 6137 3780 6141 3836
rect 6141 3780 6197 3836
rect 6197 3780 6201 3836
rect 6137 3776 6201 3780
rect 7875 3836 7939 3840
rect 7875 3780 7879 3836
rect 7879 3780 7935 3836
rect 7935 3780 7939 3836
rect 7875 3776 7939 3780
rect 7955 3836 8019 3840
rect 7955 3780 7959 3836
rect 7959 3780 8015 3836
rect 8015 3780 8019 3836
rect 7955 3776 8019 3780
rect 8035 3836 8099 3840
rect 8035 3780 8039 3836
rect 8039 3780 8095 3836
rect 8095 3780 8099 3836
rect 8035 3776 8099 3780
rect 8115 3836 8179 3840
rect 8115 3780 8119 3836
rect 8119 3780 8175 3836
rect 8175 3780 8179 3836
rect 8115 3776 8179 3780
rect 2601 3292 2665 3296
rect 2601 3236 2605 3292
rect 2605 3236 2661 3292
rect 2661 3236 2665 3292
rect 2601 3232 2665 3236
rect 2681 3292 2745 3296
rect 2681 3236 2685 3292
rect 2685 3236 2741 3292
rect 2741 3236 2745 3292
rect 2681 3232 2745 3236
rect 2761 3292 2825 3296
rect 2761 3236 2765 3292
rect 2765 3236 2821 3292
rect 2821 3236 2825 3292
rect 2761 3232 2825 3236
rect 2841 3292 2905 3296
rect 2841 3236 2845 3292
rect 2845 3236 2901 3292
rect 2901 3236 2905 3292
rect 2841 3232 2905 3236
rect 4579 3292 4643 3296
rect 4579 3236 4583 3292
rect 4583 3236 4639 3292
rect 4639 3236 4643 3292
rect 4579 3232 4643 3236
rect 4659 3292 4723 3296
rect 4659 3236 4663 3292
rect 4663 3236 4719 3292
rect 4719 3236 4723 3292
rect 4659 3232 4723 3236
rect 4739 3292 4803 3296
rect 4739 3236 4743 3292
rect 4743 3236 4799 3292
rect 4799 3236 4803 3292
rect 4739 3232 4803 3236
rect 4819 3292 4883 3296
rect 4819 3236 4823 3292
rect 4823 3236 4879 3292
rect 4879 3236 4883 3292
rect 4819 3232 4883 3236
rect 6557 3292 6621 3296
rect 6557 3236 6561 3292
rect 6561 3236 6617 3292
rect 6617 3236 6621 3292
rect 6557 3232 6621 3236
rect 6637 3292 6701 3296
rect 6637 3236 6641 3292
rect 6641 3236 6697 3292
rect 6697 3236 6701 3292
rect 6637 3232 6701 3236
rect 6717 3292 6781 3296
rect 6717 3236 6721 3292
rect 6721 3236 6777 3292
rect 6777 3236 6781 3292
rect 6717 3232 6781 3236
rect 6797 3292 6861 3296
rect 6797 3236 6801 3292
rect 6801 3236 6857 3292
rect 6857 3236 6861 3292
rect 6797 3232 6861 3236
rect 8535 3292 8599 3296
rect 8535 3236 8539 3292
rect 8539 3236 8595 3292
rect 8595 3236 8599 3292
rect 8535 3232 8599 3236
rect 8615 3292 8679 3296
rect 8615 3236 8619 3292
rect 8619 3236 8675 3292
rect 8675 3236 8679 3292
rect 8615 3232 8679 3236
rect 8695 3292 8759 3296
rect 8695 3236 8699 3292
rect 8699 3236 8755 3292
rect 8755 3236 8759 3292
rect 8695 3232 8759 3236
rect 8775 3292 8839 3296
rect 8775 3236 8779 3292
rect 8779 3236 8835 3292
rect 8835 3236 8839 3292
rect 8775 3232 8839 3236
rect 1941 2748 2005 2752
rect 1941 2692 1945 2748
rect 1945 2692 2001 2748
rect 2001 2692 2005 2748
rect 1941 2688 2005 2692
rect 2021 2748 2085 2752
rect 2021 2692 2025 2748
rect 2025 2692 2081 2748
rect 2081 2692 2085 2748
rect 2021 2688 2085 2692
rect 2101 2748 2165 2752
rect 2101 2692 2105 2748
rect 2105 2692 2161 2748
rect 2161 2692 2165 2748
rect 2101 2688 2165 2692
rect 2181 2748 2245 2752
rect 2181 2692 2185 2748
rect 2185 2692 2241 2748
rect 2241 2692 2245 2748
rect 2181 2688 2245 2692
rect 3919 2748 3983 2752
rect 3919 2692 3923 2748
rect 3923 2692 3979 2748
rect 3979 2692 3983 2748
rect 3919 2688 3983 2692
rect 3999 2748 4063 2752
rect 3999 2692 4003 2748
rect 4003 2692 4059 2748
rect 4059 2692 4063 2748
rect 3999 2688 4063 2692
rect 4079 2748 4143 2752
rect 4079 2692 4083 2748
rect 4083 2692 4139 2748
rect 4139 2692 4143 2748
rect 4079 2688 4143 2692
rect 4159 2748 4223 2752
rect 4159 2692 4163 2748
rect 4163 2692 4219 2748
rect 4219 2692 4223 2748
rect 4159 2688 4223 2692
rect 5897 2748 5961 2752
rect 5897 2692 5901 2748
rect 5901 2692 5957 2748
rect 5957 2692 5961 2748
rect 5897 2688 5961 2692
rect 5977 2748 6041 2752
rect 5977 2692 5981 2748
rect 5981 2692 6037 2748
rect 6037 2692 6041 2748
rect 5977 2688 6041 2692
rect 6057 2748 6121 2752
rect 6057 2692 6061 2748
rect 6061 2692 6117 2748
rect 6117 2692 6121 2748
rect 6057 2688 6121 2692
rect 6137 2748 6201 2752
rect 6137 2692 6141 2748
rect 6141 2692 6197 2748
rect 6197 2692 6201 2748
rect 6137 2688 6201 2692
rect 7875 2748 7939 2752
rect 7875 2692 7879 2748
rect 7879 2692 7935 2748
rect 7935 2692 7939 2748
rect 7875 2688 7939 2692
rect 7955 2748 8019 2752
rect 7955 2692 7959 2748
rect 7959 2692 8015 2748
rect 8015 2692 8019 2748
rect 7955 2688 8019 2692
rect 8035 2748 8099 2752
rect 8035 2692 8039 2748
rect 8039 2692 8095 2748
rect 8095 2692 8099 2748
rect 8035 2688 8099 2692
rect 8115 2748 8179 2752
rect 8115 2692 8119 2748
rect 8119 2692 8175 2748
rect 8175 2692 8179 2748
rect 8115 2688 8179 2692
rect 2601 2204 2665 2208
rect 2601 2148 2605 2204
rect 2605 2148 2661 2204
rect 2661 2148 2665 2204
rect 2601 2144 2665 2148
rect 2681 2204 2745 2208
rect 2681 2148 2685 2204
rect 2685 2148 2741 2204
rect 2741 2148 2745 2204
rect 2681 2144 2745 2148
rect 2761 2204 2825 2208
rect 2761 2148 2765 2204
rect 2765 2148 2821 2204
rect 2821 2148 2825 2204
rect 2761 2144 2825 2148
rect 2841 2204 2905 2208
rect 2841 2148 2845 2204
rect 2845 2148 2901 2204
rect 2901 2148 2905 2204
rect 2841 2144 2905 2148
rect 4579 2204 4643 2208
rect 4579 2148 4583 2204
rect 4583 2148 4639 2204
rect 4639 2148 4643 2204
rect 4579 2144 4643 2148
rect 4659 2204 4723 2208
rect 4659 2148 4663 2204
rect 4663 2148 4719 2204
rect 4719 2148 4723 2204
rect 4659 2144 4723 2148
rect 4739 2204 4803 2208
rect 4739 2148 4743 2204
rect 4743 2148 4799 2204
rect 4799 2148 4803 2204
rect 4739 2144 4803 2148
rect 4819 2204 4883 2208
rect 4819 2148 4823 2204
rect 4823 2148 4879 2204
rect 4879 2148 4883 2204
rect 4819 2144 4883 2148
rect 6557 2204 6621 2208
rect 6557 2148 6561 2204
rect 6561 2148 6617 2204
rect 6617 2148 6621 2204
rect 6557 2144 6621 2148
rect 6637 2204 6701 2208
rect 6637 2148 6641 2204
rect 6641 2148 6697 2204
rect 6697 2148 6701 2204
rect 6637 2144 6701 2148
rect 6717 2204 6781 2208
rect 6717 2148 6721 2204
rect 6721 2148 6777 2204
rect 6777 2148 6781 2204
rect 6717 2144 6781 2148
rect 6797 2204 6861 2208
rect 6797 2148 6801 2204
rect 6801 2148 6857 2204
rect 6857 2148 6861 2204
rect 6797 2144 6861 2148
rect 8535 2204 8599 2208
rect 8535 2148 8539 2204
rect 8539 2148 8595 2204
rect 8595 2148 8599 2204
rect 8535 2144 8599 2148
rect 8615 2204 8679 2208
rect 8615 2148 8619 2204
rect 8619 2148 8675 2204
rect 8675 2148 8679 2204
rect 8615 2144 8679 2148
rect 8695 2204 8759 2208
rect 8695 2148 8699 2204
rect 8699 2148 8755 2204
rect 8755 2148 8759 2204
rect 8695 2144 8759 2148
rect 8775 2204 8839 2208
rect 8775 2148 8779 2204
rect 8779 2148 8835 2204
rect 8835 2148 8839 2204
rect 8775 2144 8839 2148
<< metal4 >>
rect 1933 9280 2253 9840
rect 1933 9216 1941 9280
rect 2005 9216 2021 9280
rect 2085 9216 2101 9280
rect 2165 9216 2181 9280
rect 2245 9216 2253 9280
rect 1933 8958 2253 9216
rect 1933 8722 1975 8958
rect 2211 8722 2253 8958
rect 1933 8192 2253 8722
rect 1933 8128 1941 8192
rect 2005 8128 2021 8192
rect 2085 8128 2101 8192
rect 2165 8128 2181 8192
rect 2245 8128 2253 8192
rect 1933 7104 2253 8128
rect 1933 7040 1941 7104
rect 2005 7054 2021 7104
rect 2085 7054 2101 7104
rect 2165 7054 2181 7104
rect 2245 7040 2253 7104
rect 1933 6818 1975 7040
rect 2211 6818 2253 7040
rect 1933 6016 2253 6818
rect 1933 5952 1941 6016
rect 2005 5952 2021 6016
rect 2085 5952 2101 6016
rect 2165 5952 2181 6016
rect 2245 5952 2253 6016
rect 1933 5150 2253 5952
rect 1933 4928 1975 5150
rect 2211 4928 2253 5150
rect 1933 4864 1941 4928
rect 2005 4864 2021 4914
rect 2085 4864 2101 4914
rect 2165 4864 2181 4914
rect 2245 4864 2253 4928
rect 1933 3840 2253 4864
rect 1933 3776 1941 3840
rect 2005 3776 2021 3840
rect 2085 3776 2101 3840
rect 2165 3776 2181 3840
rect 2245 3776 2253 3840
rect 1933 3246 2253 3776
rect 1933 3010 1975 3246
rect 2211 3010 2253 3246
rect 1933 2752 2253 3010
rect 1933 2688 1941 2752
rect 2005 2688 2021 2752
rect 2085 2688 2101 2752
rect 2165 2688 2181 2752
rect 2245 2688 2253 2752
rect 1933 2128 2253 2688
rect 2593 9824 2913 9840
rect 2593 9760 2601 9824
rect 2665 9760 2681 9824
rect 2745 9760 2761 9824
rect 2825 9760 2841 9824
rect 2905 9760 2913 9824
rect 2593 9618 2913 9760
rect 2593 9382 2635 9618
rect 2871 9382 2913 9618
rect 2593 8736 2913 9382
rect 2593 8672 2601 8736
rect 2665 8672 2681 8736
rect 2745 8672 2761 8736
rect 2825 8672 2841 8736
rect 2905 8672 2913 8736
rect 2593 7714 2913 8672
rect 2593 7648 2635 7714
rect 2871 7648 2913 7714
rect 2593 7584 2601 7648
rect 2905 7584 2913 7648
rect 2593 7478 2635 7584
rect 2871 7478 2913 7584
rect 2593 6560 2913 7478
rect 2593 6496 2601 6560
rect 2665 6496 2681 6560
rect 2745 6496 2761 6560
rect 2825 6496 2841 6560
rect 2905 6496 2913 6560
rect 2593 5810 2913 6496
rect 2593 5574 2635 5810
rect 2871 5574 2913 5810
rect 2593 5472 2913 5574
rect 2593 5408 2601 5472
rect 2665 5408 2681 5472
rect 2745 5408 2761 5472
rect 2825 5408 2841 5472
rect 2905 5408 2913 5472
rect 2593 4384 2913 5408
rect 2593 4320 2601 4384
rect 2665 4320 2681 4384
rect 2745 4320 2761 4384
rect 2825 4320 2841 4384
rect 2905 4320 2913 4384
rect 2593 3906 2913 4320
rect 2593 3670 2635 3906
rect 2871 3670 2913 3906
rect 2593 3296 2913 3670
rect 2593 3232 2601 3296
rect 2665 3232 2681 3296
rect 2745 3232 2761 3296
rect 2825 3232 2841 3296
rect 2905 3232 2913 3296
rect 2593 2208 2913 3232
rect 2593 2144 2601 2208
rect 2665 2144 2681 2208
rect 2745 2144 2761 2208
rect 2825 2144 2841 2208
rect 2905 2144 2913 2208
rect 2593 2128 2913 2144
rect 3911 9280 4231 9840
rect 3911 9216 3919 9280
rect 3983 9216 3999 9280
rect 4063 9216 4079 9280
rect 4143 9216 4159 9280
rect 4223 9216 4231 9280
rect 3911 8958 4231 9216
rect 3911 8722 3953 8958
rect 4189 8722 4231 8958
rect 3911 8192 4231 8722
rect 3911 8128 3919 8192
rect 3983 8128 3999 8192
rect 4063 8128 4079 8192
rect 4143 8128 4159 8192
rect 4223 8128 4231 8192
rect 3911 7104 4231 8128
rect 3911 7040 3919 7104
rect 3983 7054 3999 7104
rect 4063 7054 4079 7104
rect 4143 7054 4159 7104
rect 4223 7040 4231 7104
rect 3911 6818 3953 7040
rect 4189 6818 4231 7040
rect 3911 6016 4231 6818
rect 3911 5952 3919 6016
rect 3983 5952 3999 6016
rect 4063 5952 4079 6016
rect 4143 5952 4159 6016
rect 4223 5952 4231 6016
rect 3911 5150 4231 5952
rect 3911 4928 3953 5150
rect 4189 4928 4231 5150
rect 3911 4864 3919 4928
rect 3983 4864 3999 4914
rect 4063 4864 4079 4914
rect 4143 4864 4159 4914
rect 4223 4864 4231 4928
rect 3911 3840 4231 4864
rect 3911 3776 3919 3840
rect 3983 3776 3999 3840
rect 4063 3776 4079 3840
rect 4143 3776 4159 3840
rect 4223 3776 4231 3840
rect 3911 3246 4231 3776
rect 3911 3010 3953 3246
rect 4189 3010 4231 3246
rect 3911 2752 4231 3010
rect 3911 2688 3919 2752
rect 3983 2688 3999 2752
rect 4063 2688 4079 2752
rect 4143 2688 4159 2752
rect 4223 2688 4231 2752
rect 3911 2128 4231 2688
rect 4571 9824 4891 9840
rect 4571 9760 4579 9824
rect 4643 9760 4659 9824
rect 4723 9760 4739 9824
rect 4803 9760 4819 9824
rect 4883 9760 4891 9824
rect 4571 9618 4891 9760
rect 4571 9382 4613 9618
rect 4849 9382 4891 9618
rect 4571 8736 4891 9382
rect 4571 8672 4579 8736
rect 4643 8672 4659 8736
rect 4723 8672 4739 8736
rect 4803 8672 4819 8736
rect 4883 8672 4891 8736
rect 4571 7714 4891 8672
rect 4571 7648 4613 7714
rect 4849 7648 4891 7714
rect 4571 7584 4579 7648
rect 4883 7584 4891 7648
rect 4571 7478 4613 7584
rect 4849 7478 4891 7584
rect 4571 6560 4891 7478
rect 4571 6496 4579 6560
rect 4643 6496 4659 6560
rect 4723 6496 4739 6560
rect 4803 6496 4819 6560
rect 4883 6496 4891 6560
rect 4571 5810 4891 6496
rect 4571 5574 4613 5810
rect 4849 5574 4891 5810
rect 4571 5472 4891 5574
rect 4571 5408 4579 5472
rect 4643 5408 4659 5472
rect 4723 5408 4739 5472
rect 4803 5408 4819 5472
rect 4883 5408 4891 5472
rect 4571 4384 4891 5408
rect 4571 4320 4579 4384
rect 4643 4320 4659 4384
rect 4723 4320 4739 4384
rect 4803 4320 4819 4384
rect 4883 4320 4891 4384
rect 4571 3906 4891 4320
rect 4571 3670 4613 3906
rect 4849 3670 4891 3906
rect 4571 3296 4891 3670
rect 4571 3232 4579 3296
rect 4643 3232 4659 3296
rect 4723 3232 4739 3296
rect 4803 3232 4819 3296
rect 4883 3232 4891 3296
rect 4571 2208 4891 3232
rect 4571 2144 4579 2208
rect 4643 2144 4659 2208
rect 4723 2144 4739 2208
rect 4803 2144 4819 2208
rect 4883 2144 4891 2208
rect 4571 2128 4891 2144
rect 5889 9280 6209 9840
rect 5889 9216 5897 9280
rect 5961 9216 5977 9280
rect 6041 9216 6057 9280
rect 6121 9216 6137 9280
rect 6201 9216 6209 9280
rect 5889 8958 6209 9216
rect 5889 8722 5931 8958
rect 6167 8722 6209 8958
rect 5889 8192 6209 8722
rect 5889 8128 5897 8192
rect 5961 8128 5977 8192
rect 6041 8128 6057 8192
rect 6121 8128 6137 8192
rect 6201 8128 6209 8192
rect 5889 7104 6209 8128
rect 5889 7040 5897 7104
rect 5961 7054 5977 7104
rect 6041 7054 6057 7104
rect 6121 7054 6137 7104
rect 6201 7040 6209 7104
rect 5889 6818 5931 7040
rect 6167 6818 6209 7040
rect 5889 6016 6209 6818
rect 5889 5952 5897 6016
rect 5961 5952 5977 6016
rect 6041 5952 6057 6016
rect 6121 5952 6137 6016
rect 6201 5952 6209 6016
rect 5889 5150 6209 5952
rect 5889 4928 5931 5150
rect 6167 4928 6209 5150
rect 5889 4864 5897 4928
rect 5961 4864 5977 4914
rect 6041 4864 6057 4914
rect 6121 4864 6137 4914
rect 6201 4864 6209 4928
rect 5889 3840 6209 4864
rect 5889 3776 5897 3840
rect 5961 3776 5977 3840
rect 6041 3776 6057 3840
rect 6121 3776 6137 3840
rect 6201 3776 6209 3840
rect 5889 3246 6209 3776
rect 5889 3010 5931 3246
rect 6167 3010 6209 3246
rect 5889 2752 6209 3010
rect 5889 2688 5897 2752
rect 5961 2688 5977 2752
rect 6041 2688 6057 2752
rect 6121 2688 6137 2752
rect 6201 2688 6209 2752
rect 5889 2128 6209 2688
rect 6549 9824 6869 9840
rect 6549 9760 6557 9824
rect 6621 9760 6637 9824
rect 6701 9760 6717 9824
rect 6781 9760 6797 9824
rect 6861 9760 6869 9824
rect 6549 9618 6869 9760
rect 6549 9382 6591 9618
rect 6827 9382 6869 9618
rect 6549 8736 6869 9382
rect 6549 8672 6557 8736
rect 6621 8672 6637 8736
rect 6701 8672 6717 8736
rect 6781 8672 6797 8736
rect 6861 8672 6869 8736
rect 6549 7714 6869 8672
rect 6549 7648 6591 7714
rect 6827 7648 6869 7714
rect 6549 7584 6557 7648
rect 6861 7584 6869 7648
rect 6549 7478 6591 7584
rect 6827 7478 6869 7584
rect 6549 6560 6869 7478
rect 6549 6496 6557 6560
rect 6621 6496 6637 6560
rect 6701 6496 6717 6560
rect 6781 6496 6797 6560
rect 6861 6496 6869 6560
rect 6549 5810 6869 6496
rect 6549 5574 6591 5810
rect 6827 5574 6869 5810
rect 6549 5472 6869 5574
rect 6549 5408 6557 5472
rect 6621 5408 6637 5472
rect 6701 5408 6717 5472
rect 6781 5408 6797 5472
rect 6861 5408 6869 5472
rect 6549 4384 6869 5408
rect 6549 4320 6557 4384
rect 6621 4320 6637 4384
rect 6701 4320 6717 4384
rect 6781 4320 6797 4384
rect 6861 4320 6869 4384
rect 6549 3906 6869 4320
rect 6549 3670 6591 3906
rect 6827 3670 6869 3906
rect 6549 3296 6869 3670
rect 6549 3232 6557 3296
rect 6621 3232 6637 3296
rect 6701 3232 6717 3296
rect 6781 3232 6797 3296
rect 6861 3232 6869 3296
rect 6549 2208 6869 3232
rect 6549 2144 6557 2208
rect 6621 2144 6637 2208
rect 6701 2144 6717 2208
rect 6781 2144 6797 2208
rect 6861 2144 6869 2208
rect 6549 2128 6869 2144
rect 7867 9280 8187 9840
rect 7867 9216 7875 9280
rect 7939 9216 7955 9280
rect 8019 9216 8035 9280
rect 8099 9216 8115 9280
rect 8179 9216 8187 9280
rect 7867 8958 8187 9216
rect 7867 8722 7909 8958
rect 8145 8722 8187 8958
rect 7867 8192 8187 8722
rect 7867 8128 7875 8192
rect 7939 8128 7955 8192
rect 8019 8128 8035 8192
rect 8099 8128 8115 8192
rect 8179 8128 8187 8192
rect 7867 7104 8187 8128
rect 7867 7040 7875 7104
rect 7939 7054 7955 7104
rect 8019 7054 8035 7104
rect 8099 7054 8115 7104
rect 8179 7040 8187 7104
rect 7867 6818 7909 7040
rect 8145 6818 8187 7040
rect 7867 6016 8187 6818
rect 7867 5952 7875 6016
rect 7939 5952 7955 6016
rect 8019 5952 8035 6016
rect 8099 5952 8115 6016
rect 8179 5952 8187 6016
rect 7867 5150 8187 5952
rect 7867 4928 7909 5150
rect 8145 4928 8187 5150
rect 7867 4864 7875 4928
rect 7939 4864 7955 4914
rect 8019 4864 8035 4914
rect 8099 4864 8115 4914
rect 8179 4864 8187 4928
rect 7867 3840 8187 4864
rect 7867 3776 7875 3840
rect 7939 3776 7955 3840
rect 8019 3776 8035 3840
rect 8099 3776 8115 3840
rect 8179 3776 8187 3840
rect 7867 3246 8187 3776
rect 7867 3010 7909 3246
rect 8145 3010 8187 3246
rect 7867 2752 8187 3010
rect 7867 2688 7875 2752
rect 7939 2688 7955 2752
rect 8019 2688 8035 2752
rect 8099 2688 8115 2752
rect 8179 2688 8187 2752
rect 7867 2128 8187 2688
rect 8527 9824 8847 9840
rect 8527 9760 8535 9824
rect 8599 9760 8615 9824
rect 8679 9760 8695 9824
rect 8759 9760 8775 9824
rect 8839 9760 8847 9824
rect 8527 9618 8847 9760
rect 8527 9382 8569 9618
rect 8805 9382 8847 9618
rect 8527 8736 8847 9382
rect 8527 8672 8535 8736
rect 8599 8672 8615 8736
rect 8679 8672 8695 8736
rect 8759 8672 8775 8736
rect 8839 8672 8847 8736
rect 8527 7714 8847 8672
rect 8527 7648 8569 7714
rect 8805 7648 8847 7714
rect 8527 7584 8535 7648
rect 8839 7584 8847 7648
rect 8527 7478 8569 7584
rect 8805 7478 8847 7584
rect 8527 6560 8847 7478
rect 8527 6496 8535 6560
rect 8599 6496 8615 6560
rect 8679 6496 8695 6560
rect 8759 6496 8775 6560
rect 8839 6496 8847 6560
rect 8527 5810 8847 6496
rect 8527 5574 8569 5810
rect 8805 5574 8847 5810
rect 8527 5472 8847 5574
rect 8527 5408 8535 5472
rect 8599 5408 8615 5472
rect 8679 5408 8695 5472
rect 8759 5408 8775 5472
rect 8839 5408 8847 5472
rect 8527 4384 8847 5408
rect 8527 4320 8535 4384
rect 8599 4320 8615 4384
rect 8679 4320 8695 4384
rect 8759 4320 8775 4384
rect 8839 4320 8847 4384
rect 8527 3906 8847 4320
rect 8527 3670 8569 3906
rect 8805 3670 8847 3906
rect 8527 3296 8847 3670
rect 8527 3232 8535 3296
rect 8599 3232 8615 3296
rect 8679 3232 8695 3296
rect 8759 3232 8775 3296
rect 8839 3232 8847 3296
rect 8527 2208 8847 3232
rect 8527 2144 8535 2208
rect 8599 2144 8615 2208
rect 8679 2144 8695 2208
rect 8759 2144 8775 2208
rect 8839 2144 8847 2208
rect 8527 2128 8847 2144
<< via4 >>
rect 1975 8722 2211 8958
rect 1975 7040 2005 7054
rect 2005 7040 2021 7054
rect 2021 7040 2085 7054
rect 2085 7040 2101 7054
rect 2101 7040 2165 7054
rect 2165 7040 2181 7054
rect 2181 7040 2211 7054
rect 1975 6818 2211 7040
rect 1975 4928 2211 5150
rect 1975 4914 2005 4928
rect 2005 4914 2021 4928
rect 2021 4914 2085 4928
rect 2085 4914 2101 4928
rect 2101 4914 2165 4928
rect 2165 4914 2181 4928
rect 2181 4914 2211 4928
rect 1975 3010 2211 3246
rect 2635 9382 2871 9618
rect 2635 7648 2871 7714
rect 2635 7584 2665 7648
rect 2665 7584 2681 7648
rect 2681 7584 2745 7648
rect 2745 7584 2761 7648
rect 2761 7584 2825 7648
rect 2825 7584 2841 7648
rect 2841 7584 2871 7648
rect 2635 7478 2871 7584
rect 2635 5574 2871 5810
rect 2635 3670 2871 3906
rect 3953 8722 4189 8958
rect 3953 7040 3983 7054
rect 3983 7040 3999 7054
rect 3999 7040 4063 7054
rect 4063 7040 4079 7054
rect 4079 7040 4143 7054
rect 4143 7040 4159 7054
rect 4159 7040 4189 7054
rect 3953 6818 4189 7040
rect 3953 4928 4189 5150
rect 3953 4914 3983 4928
rect 3983 4914 3999 4928
rect 3999 4914 4063 4928
rect 4063 4914 4079 4928
rect 4079 4914 4143 4928
rect 4143 4914 4159 4928
rect 4159 4914 4189 4928
rect 3953 3010 4189 3246
rect 4613 9382 4849 9618
rect 4613 7648 4849 7714
rect 4613 7584 4643 7648
rect 4643 7584 4659 7648
rect 4659 7584 4723 7648
rect 4723 7584 4739 7648
rect 4739 7584 4803 7648
rect 4803 7584 4819 7648
rect 4819 7584 4849 7648
rect 4613 7478 4849 7584
rect 4613 5574 4849 5810
rect 4613 3670 4849 3906
rect 5931 8722 6167 8958
rect 5931 7040 5961 7054
rect 5961 7040 5977 7054
rect 5977 7040 6041 7054
rect 6041 7040 6057 7054
rect 6057 7040 6121 7054
rect 6121 7040 6137 7054
rect 6137 7040 6167 7054
rect 5931 6818 6167 7040
rect 5931 4928 6167 5150
rect 5931 4914 5961 4928
rect 5961 4914 5977 4928
rect 5977 4914 6041 4928
rect 6041 4914 6057 4928
rect 6057 4914 6121 4928
rect 6121 4914 6137 4928
rect 6137 4914 6167 4928
rect 5931 3010 6167 3246
rect 6591 9382 6827 9618
rect 6591 7648 6827 7714
rect 6591 7584 6621 7648
rect 6621 7584 6637 7648
rect 6637 7584 6701 7648
rect 6701 7584 6717 7648
rect 6717 7584 6781 7648
rect 6781 7584 6797 7648
rect 6797 7584 6827 7648
rect 6591 7478 6827 7584
rect 6591 5574 6827 5810
rect 6591 3670 6827 3906
rect 7909 8722 8145 8958
rect 7909 7040 7939 7054
rect 7939 7040 7955 7054
rect 7955 7040 8019 7054
rect 8019 7040 8035 7054
rect 8035 7040 8099 7054
rect 8099 7040 8115 7054
rect 8115 7040 8145 7054
rect 7909 6818 8145 7040
rect 7909 4928 8145 5150
rect 7909 4914 7939 4928
rect 7939 4914 7955 4928
rect 7955 4914 8019 4928
rect 8019 4914 8035 4928
rect 8035 4914 8099 4928
rect 8099 4914 8115 4928
rect 8115 4914 8145 4928
rect 7909 3010 8145 3246
rect 8569 9382 8805 9618
rect 8569 7648 8805 7714
rect 8569 7584 8599 7648
rect 8599 7584 8615 7648
rect 8615 7584 8679 7648
rect 8679 7584 8695 7648
rect 8695 7584 8759 7648
rect 8759 7584 8775 7648
rect 8775 7584 8805 7648
rect 8569 7478 8805 7584
rect 8569 5574 8805 5810
rect 8569 3670 8805 3906
<< metal5 >>
rect 1056 9618 9064 9660
rect 1056 9382 2635 9618
rect 2871 9382 4613 9618
rect 4849 9382 6591 9618
rect 6827 9382 8569 9618
rect 8805 9382 9064 9618
rect 1056 9340 9064 9382
rect 1056 8958 9064 9000
rect 1056 8722 1975 8958
rect 2211 8722 3953 8958
rect 4189 8722 5931 8958
rect 6167 8722 7909 8958
rect 8145 8722 9064 8958
rect 1056 8680 9064 8722
rect 1056 7714 9064 7756
rect 1056 7478 2635 7714
rect 2871 7478 4613 7714
rect 4849 7478 6591 7714
rect 6827 7478 8569 7714
rect 8805 7478 9064 7714
rect 1056 7436 9064 7478
rect 1056 7054 9064 7096
rect 1056 6818 1975 7054
rect 2211 6818 3953 7054
rect 4189 6818 5931 7054
rect 6167 6818 7909 7054
rect 8145 6818 9064 7054
rect 1056 6776 9064 6818
rect 1056 5810 9064 5852
rect 1056 5574 2635 5810
rect 2871 5574 4613 5810
rect 4849 5574 6591 5810
rect 6827 5574 8569 5810
rect 8805 5574 9064 5810
rect 1056 5532 9064 5574
rect 1056 5150 9064 5192
rect 1056 4914 1975 5150
rect 2211 4914 3953 5150
rect 4189 4914 5931 5150
rect 6167 4914 7909 5150
rect 8145 4914 9064 5150
rect 1056 4872 9064 4914
rect 1056 3906 9064 3948
rect 1056 3670 2635 3906
rect 2871 3670 4613 3906
rect 4849 3670 6591 3906
rect 6827 3670 8569 3906
rect 8805 3670 9064 3906
rect 1056 3628 9064 3670
rect 1056 3246 9064 3288
rect 1056 3010 1975 3246
rect 2211 3010 3953 3246
rect 4189 3010 5931 3246
rect 6167 3010 7909 3246
rect 8145 3010 9064 3246
rect 1056 2968 9064 3010
use sky130_fd_sc_hd__clkbuf_4  _092_ ASIC/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 7544 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _093_ ASIC/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 7268 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__nand3_4  _094_ ASIC/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 5796 0 -1 4352
box -38 -48 1326 592
use sky130_fd_sc_hd__o2111a_1  _095_ ASIC/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 5060 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _096_ ASIC/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5152 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _097_ ASIC/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 5612 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _098_ ASIC/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 6348 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _099_ ASIC/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 2668 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__nand4_4  _100_ ASIC/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 5336 0 1 6528
box -38 -48 1602 592
use sky130_fd_sc_hd__a22oi_4  _101_ ASIC/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5612 0 1 6528
box -38 -48 1602 592
use sky130_fd_sc_hd__and3b_1  _102_ ASIC/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 5612 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _103_ ASIC/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 7452 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _104_ ASIC/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 2300 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _105_ ASIC/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 6440 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _106_ ASIC/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 6348 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _107_
timestamp 1688980957
transform 1 0 8372 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__nand4b_2  _108_ ASIC/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 8004 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__o211a_1  _109_ ASIC/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 6256 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _110_ ASIC/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 7912 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__nand4_1  _111_ ASIC/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3772 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__a2bb2oi_1  _112_ ASIC/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 6992 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _113_
timestamp 1688980957
transform 1 0 5796 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _114_ ASIC/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 8648 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a31oi_1  _115_ ASIC/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 8372 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _116_ ASIC/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 1748 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _117_ ASIC/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 6808 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__or2b_1  _118_ ASIC/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 6440 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _119_
timestamp 1688980957
transform -1 0 4324 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _120_
timestamp 1688980957
transform 1 0 4324 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _121_
timestamp 1688980957
transform -1 0 8740 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nand3b_1  _122_ ASIC/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 8648 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__nand4_1  _123_
timestamp 1688980957
transform 1 0 5704 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _124_
timestamp 1688980957
transform 1 0 3404 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__o311a_1  _125_ ASIC/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5336 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _126_
timestamp 1688980957
transform 1 0 5060 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _127_
timestamp 1688980957
transform 1 0 3312 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__o21bai_1  _128_ ASIC/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 6808 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _129_
timestamp 1688980957
transform 1 0 3956 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a32oi_1  _130_ ASIC/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5612 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__o2111ai_1  _131_ ASIC/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4232 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a22oi_1  _132_ ASIC/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 3404 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_2  _133_ ASIC/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5244 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _134_ ASIC/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 6256 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _135_ ASIC/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 7452 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a41oi_2  _136_ ASIC/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 4416 0 -1 6528
box -38 -48 1234 592
use sky130_fd_sc_hd__or2_1  _137_
timestamp 1688980957
transform 1 0 4968 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _138_
timestamp 1688980957
transform -1 0 6716 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _139_
timestamp 1688980957
transform 1 0 5704 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _140_
timestamp 1688980957
transform -1 0 3680 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _141_ ASIC/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 6348 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _142_ ASIC/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3772 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _143_
timestamp 1688980957
transform -1 0 2484 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__nand4_2  _144_ ASIC/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 2392 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__a32o_1  _145_
timestamp 1688980957
transform 1 0 2944 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _146_ ASIC/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1380 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a41o_1  _147_ ASIC/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 2852 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _148_
timestamp 1688980957
transform 1 0 1932 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__nor3_1  _149_ ASIC/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3312 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _150_
timestamp 1688980957
transform 1 0 2208 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _151_
timestamp 1688980957
transform 1 0 1380 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _152_ ASIC/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1564 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_2  _153_ ASIC/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3496 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _154_
timestamp 1688980957
transform 1 0 4600 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a31oi_1  _155_
timestamp 1688980957
transform -1 0 3312 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__o211ai_2  _156_ ASIC/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3772 0 1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__o2111ai_1  _157_
timestamp 1688980957
transform 1 0 1932 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a22oi_1  _158_
timestamp 1688980957
transform -1 0 2576 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _159_ ASIC/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 5244 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _160_ ASIC/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1564 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__a32oi_1  _161_
timestamp 1688980957
transform 1 0 2852 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a211oi_2  _162_ ASIC/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 7268 0 -1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__a31oi_1  _163_
timestamp 1688980957
transform 1 0 6532 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _164_
timestamp 1688980957
transform 1 0 7820 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _165_
timestamp 1688980957
transform 1 0 8464 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _166_
timestamp 1688980957
transform 1 0 8188 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__o2111ai_1  _167_
timestamp 1688980957
transform 1 0 6808 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _168_ ASIC/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 7820 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__and3b_1  _169_
timestamp 1688980957
transform -1 0 8464 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _170_
timestamp 1688980957
transform -1 0 8740 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _171_
timestamp 1688980957
transform 1 0 8372 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__o2111a_1  _172_
timestamp 1688980957
transform 1 0 6992 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__o2bb2ai_1  _173_ ASIC/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 7176 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _174_
timestamp 1688980957
transform -1 0 2024 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_4  _175_ ASIC/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 5704 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_4  _176_ ASIC/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1380 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _177_
timestamp 1688980957
transform -1 0 2208 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_4  _178_
timestamp 1688980957
transform 1 0 4416 0 -1 7616
box -38 -48 1326 592
use sky130_fd_sc_hd__and2b_2  _179_ ASIC/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 6348 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_4  _180_ ASIC/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4140 0 -1 5440
box -38 -48 1234 592
use sky130_fd_sc_hd__clkbuf_4  _181_
timestamp 1688980957
transform 1 0 6992 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _182_
timestamp 1688980957
transform 1 0 7544 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_2  _183_ ASIC/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 4508 0 -1 4352
box -38 -48 1234 592
use sky130_fd_sc_hd__dfxtp_2  _184_ ASIC/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 5336 0 1 2176
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _185_ ASIC/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 7268 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _186_
timestamp 1688980957
transform 1 0 5336 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _187_
timestamp 1688980957
transform 1 0 6992 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _188_
timestamp 1688980957
transform -1 0 2852 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_4  _189_ ASIC/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 7452 0 1 8704
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_2  _190_
timestamp 1688980957
transform -1 0 5704 0 1 8704
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _191_
timestamp 1688980957
transform 1 0 3312 0 -1 8704
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _192_
timestamp 1688980957
transform -1 0 2944 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _193_
timestamp 1688980957
transform -1 0 2852 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _194_
timestamp 1688980957
transform 1 0 1380 0 1 6528
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _195_
timestamp 1688980957
transform 1 0 1380 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _196_
timestamp 1688980957
transform 1 0 1380 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _197_
timestamp 1688980957
transform 1 0 7268 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _198_
timestamp 1688980957
transform 1 0 7268 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _199_
timestamp 1688980957
transform 1 0 7268 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk ASIC/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4416 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_clk
timestamp 1688980957
transform -1 0 4416 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_clk
timestamp 1688980957
transform -1 0 4416 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_46 ASIC/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5336 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_82 ASIC/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 8648 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_9
timestamp 1688980957
transform 1 0 1932 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_57
timestamp 1688980957
transform 1 0 6348 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_82
timestamp 1688980957
transform 1 0 8648 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_3
timestamp 1688980957
transform 1 0 1380 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_3
timestamp 1688980957
transform 1 0 1380 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_29
timestamp 1688980957
transform 1 0 3772 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_41
timestamp 1688980957
transform 1 0 4876 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_70
timestamp 1688980957
transform 1 0 7544 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_79
timestamp 1688980957
transform 1 0 8372 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_54
timestamp 1688980957
transform 1 0 6072 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_78
timestamp 1688980957
transform 1 0 8280 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_3
timestamp 1688980957
transform 1 0 1380 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_11
timestamp 1688980957
transform 1 0 2116 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_26
timestamp 1688980957
transform 1 0 3496 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_58
timestamp 1688980957
transform 1 0 6440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_73
timestamp 1688980957
transform 1 0 7820 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_16
timestamp 1688980957
transform 1 0 2576 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_12
timestamp 1688980957
transform 1 0 2208 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_55
timestamp 1688980957
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_82
timestamp 1688980957
transform 1 0 8648 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 1688980957
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_61
timestamp 1688980957
transform 1 0 6716 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_81
timestamp 1688980957
transform 1 0 8556 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_12
timestamp 1688980957
transform 1 0 2208 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_41
timestamp 1688980957
transform 1 0 4876 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_65
timestamp 1688980957
transform 1 0 7084 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_3
timestamp 1688980957
transform 1 0 1380 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_29 ASIC/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3772 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_3
timestamp 1688980957
transform 1 0 1380 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_23
timestamp 1688980957
transform 1 0 3220 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_40 ASIC/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4784 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_51
timestamp 1688980957
transform 1 0 5796 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_55
timestamp 1688980957
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_65
timestamp 1688980957
transform 1 0 7084 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8 ASIC/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 3496 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 1688980957
transform -1 0 8740 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold10
timestamp 1688980957
transform -1 0 5152 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp 1688980957
transform 1 0 5520 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold13
timestamp 1688980957
transform -1 0 8372 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold14
timestamp 1688980957
transform -1 0 3312 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold16
timestamp 1688980957
transform 1 0 7728 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold17
timestamp 1688980957
transform -1 0 7084 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold18
timestamp 1688980957
transform -1 0 3680 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold19
timestamp 1688980957
transform 1 0 2484 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold20
timestamp 1688980957
transform -1 0 8280 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold24
timestamp 1688980957
transform -1 0 3312 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  input1 ASIC/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 8740 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input2
timestamp 1688980957
transform 1 0 6808 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input3
timestamp 1688980957
transform 1 0 2024 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  output4
timestamp 1688980957
transform -1 0 1932 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_0 ASIC/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1688980957
transform -1 0 9016 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1688980957
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1688980957
transform -1 0 9016 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1688980957
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1688980957
transform -1 0 9016 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1688980957
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1688980957
transform -1 0 9016 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1688980957
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1688980957
transform -1 0 9016 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1688980957
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1688980957
transform -1 0 9016 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1688980957
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1688980957
transform -1 0 9016 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1688980957
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1688980957
transform -1 0 9016 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1688980957
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1688980957
transform -1 0 9016 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1688980957
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1688980957
transform -1 0 9016 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1688980957
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1688980957
transform -1 0 9016 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1688980957
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1688980957
transform -1 0 9016 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1688980957
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1688980957
transform -1 0 9016 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1688980957
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1688980957
transform -1 0 9016 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  rebuffer1
timestamp 1688980957
transform -1 0 5796 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  rebuffer2
timestamp 1688980957
transform -1 0 4048 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  rebuffer3
timestamp 1688980957
transform -1 0 2576 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  rebuffer4
timestamp 1688980957
transform 1 0 5888 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  rebuffer5
timestamp 1688980957
transform -1 0 1840 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  rebuffer6
timestamp 1688980957
transform -1 0 4784 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_28 ASIC/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_29
timestamp 1688980957
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_30
timestamp 1688980957
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_31
timestamp 1688980957
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_32
timestamp 1688980957
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_33
timestamp 1688980957
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_34
timestamp 1688980957
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_35
timestamp 1688980957
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_36
timestamp 1688980957
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_37
timestamp 1688980957
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_38
timestamp 1688980957
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_39
timestamp 1688980957
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_40
timestamp 1688980957
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_41
timestamp 1688980957
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_42
timestamp 1688980957
transform 1 0 3680 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_43
timestamp 1688980957
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
<< labels >>
flabel metal4 s 2593 2128 2913 9840 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 4571 2128 4891 9840 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 6549 2128 6869 9840 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 8527 2128 8847 9840 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 3628 9064 3948 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 5532 9064 5852 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 7436 9064 7756 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 9340 9064 9660 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 1933 2128 2253 9840 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 3911 2128 4231 9840 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 5889 2128 6209 9840 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 7867 2128 8187 9840 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 2968 9064 3288 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 4872 9064 5192 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 6776 9064 7096 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 8680 9064 9000 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal3 s 0 8848 800 8968 0 FreeSans 480 0 0 0 clk
port 2 nsew signal input
flabel metal2 s 18 0 74 800 0 FreeSans 224 90 0 0 clkout
port 3 nsew signal tristate
flabel metal3 s 9412 7488 10212 7608 0 FreeSans 480 0 0 0 reset
port 4 nsew signal input
flabel metal2 s 5814 11556 5870 12356 0 FreeSans 224 90 0 0 sel[0]
port 5 nsew signal input
flabel metal2 s 8390 0 8446 800 0 FreeSans 224 90 0 0 sel[1]
port 6 nsew signal input
rlabel metal1 5060 9792 5060 9792 0 VGND
rlabel metal1 5060 9248 5060 9248 0 VPWR
rlabel metal1 5121 2346 5121 2346 0 _000_
rlabel metal1 7488 3502 7488 3502 0 _001_
rlabel metal1 6486 2618 6486 2618 0 _002_
rlabel metal1 7212 4114 7212 4114 0 _003_
rlabel metal1 2724 2414 2724 2414 0 _004_
rlabel metal1 7222 8942 7222 8942 0 _005_
rlabel metal2 5750 8466 5750 8466 0 _006_
rlabel metal1 3532 8466 3532 8466 0 _007_
rlabel metal1 2821 8874 2821 8874 0 _008_
rlabel metal2 2530 7106 2530 7106 0 _009_
rlabel metal1 1656 5882 1656 5882 0 _010_
rlabel metal1 2111 3502 2111 3502 0 _011_
rlabel metal1 2438 5134 2438 5134 0 _012_
rlabel via1 7585 8466 7585 8466 0 _013_
rlabel metal2 7498 8211 7498 8211 0 _014_
rlabel metal1 7534 6290 7534 6290 0 _015_
rlabel metal1 1794 6358 1794 6358 0 _016_
rlabel metal1 2116 6290 2116 6290 0 _017_
rlabel metal2 3358 5270 3358 5270 0 _018_
rlabel metal1 2024 5882 2024 5882 0 _019_
rlabel metal1 1610 5678 1610 5678 0 _020_
rlabel metal1 3450 5338 3450 5338 0 _021_
rlabel metal1 3542 4114 3542 4114 0 _022_
rlabel metal1 2162 4041 2162 4041 0 _023_
rlabel metal1 2070 4556 2070 4556 0 _024_
rlabel metal1 2162 4182 2162 4182 0 _025_
rlabel metal1 3358 5134 3358 5134 0 _026_
rlabel metal1 2484 4794 2484 4794 0 _027_
rlabel metal1 7498 6766 7498 6766 0 _028_
rlabel metal1 7268 5814 7268 5814 0 _029_
rlabel viali 7774 7855 7774 7855 0 _030_
rlabel metal1 7176 7854 7176 7854 0 _031_
rlabel metal1 7314 7922 7314 7922 0 _032_
rlabel metal1 7774 5814 7774 5814 0 _033_
rlabel metal2 8418 4726 8418 4726 0 _034_
rlabel metal1 8050 5066 8050 5066 0 _035_
rlabel metal2 7038 6256 7038 6256 0 _036_
rlabel metal2 1886 3536 1886 3536 0 _037_
rlabel metal1 4462 5134 4462 5134 0 _038_
rlabel metal1 3174 6290 3174 6290 0 _039_
rlabel metal2 4554 7038 4554 7038 0 _040_
rlabel metal1 4784 5202 4784 5202 0 _041_
rlabel metal1 6072 6290 6072 6290 0 _042_
rlabel metal2 5014 4590 5014 4590 0 _043_
rlabel metal1 5888 7378 5888 7378 0 _044_
rlabel metal1 7222 6154 7222 6154 0 _045_
rlabel metal2 4554 3774 4554 3774 0 _046_
rlabel via1 6854 7395 6854 7395 0 _047_
rlabel metal1 5520 4114 5520 4114 0 _048_
rlabel metal1 5474 3094 5474 3094 0 _049_
rlabel metal1 5106 3094 5106 3094 0 _050_
rlabel metal2 5198 5797 5198 5797 0 _051_
rlabel metal2 6946 8126 6946 8126 0 _052_
rlabel metal1 4002 6256 4002 6256 0 _053_
rlabel viali 3624 3502 3624 3502 0 _054_
rlabel metal1 7130 6766 7130 6766 0 _055_
rlabel metal1 5566 2346 5566 2346 0 _056_
rlabel metal1 6854 2890 6854 2890 0 _057_
rlabel metal2 5842 2652 5842 2652 0 _058_
rlabel metal1 6900 3162 6900 3162 0 _059_
rlabel metal1 6310 2414 6310 2414 0 _060_
rlabel metal1 5704 2414 5704 2414 0 _061_
rlabel metal1 6946 2380 6946 2380 0 _062_
rlabel metal2 7498 2006 7498 2006 0 _063_
rlabel metal2 6486 2074 6486 2074 0 _064_
rlabel metal1 6670 4250 6670 4250 0 _065_
rlabel metal2 1518 3791 1518 3791 0 _066_
rlabel metal1 1610 1836 1610 1836 0 _067_
rlabel via2 1794 3995 1794 3995 0 _068_
rlabel metal2 5658 5372 5658 5372 0 _069_
rlabel metal1 2852 5746 2852 5746 0 _070_
rlabel metal1 4738 4590 4738 4590 0 _071_
rlabel metal2 4600 4590 4600 4590 0 _072_
rlabel metal1 6853 7514 6853 7514 0 _073_
rlabel metal1 6348 7174 6348 7174 0 _074_
rlabel metal2 3542 2108 3542 2108 0 _075_
rlabel metal1 4232 2006 4232 2006 0 _076_
rlabel metal1 3634 3434 3634 3434 0 _077_
rlabel metal1 3125 2414 3125 2414 0 _078_
rlabel metal2 6486 5015 6486 5015 0 _079_
rlabel metal2 6026 4505 6026 4505 0 _080_
rlabel metal1 5750 4760 5750 4760 0 _081_
rlabel metal1 3358 2346 3358 2346 0 _082_
rlabel metal2 2346 6086 2346 6086 0 _083_
rlabel metal1 6946 8602 6946 8602 0 _084_
rlabel metal1 5014 6290 5014 6290 0 _085_
rlabel metal2 6026 7922 6026 7922 0 _086_
rlabel metal1 5934 7888 5934 7888 0 _087_
rlabel metal1 4002 9452 4002 9452 0 _088_
rlabel metal1 6021 7242 6021 7242 0 _089_
rlabel metal2 2714 9520 2714 9520 0 _090_
rlabel metal1 2576 5678 2576 5678 0 _091_
rlabel metal2 3634 7633 3634 7633 0 clk
rlabel metal2 4370 5236 4370 5236 0 clknet_0_clk
rlabel metal2 1426 4352 1426 4352 0 clknet_1_0__leaf_clk
rlabel metal2 7314 7344 7314 7344 0 clknet_1_1__leaf_clk
rlabel metal1 782 2822 782 2822 0 clkout
rlabel metal1 4370 9554 4370 9554 0 cnt1\[0\]
rlabel metal1 3404 7718 3404 7718 0 cnt1\[1\]
rlabel metal1 5014 8262 5014 8262 0 cnt1\[2\]
rlabel metal1 2806 8466 2806 8466 0 cnt1\[3\]
rlabel metal1 2116 7378 2116 7378 0 cnt1\[4\]
rlabel metal2 4646 7072 4646 7072 0 cnt1\[5\]
rlabel metal1 4600 7854 4600 7854 0 cnt2\[0\]
rlabel metal1 5106 5729 5106 5729 0 cnt2\[1\]
rlabel metal1 8326 5338 8326 5338 0 cnt3\[0\]
rlabel metal1 8510 7344 8510 7344 0 cnt3\[1\]
rlabel metal1 8832 6086 8832 6086 0 cnt3\[2\]
rlabel metal1 3772 2618 3772 2618 0 cnt4\[0\]
rlabel metal1 2346 2958 2346 2958 0 cnt4\[1\]
rlabel metal1 8464 2414 8464 2414 0 cnt4\[2\]
rlabel metal2 7866 2516 7866 2516 0 cnt4\[3\]
rlabel metal1 6394 5100 6394 5100 0 net1
rlabel metal2 6762 7140 6762 7140 0 net10
rlabel metal1 2944 5202 2944 5202 0 net12
rlabel metal1 8142 5882 8142 5882 0 net13
rlabel metal2 2622 2873 2622 2873 0 net14
rlabel metal1 6302 2822 6302 2822 0 net15
rlabel metal1 7590 4590 7590 4590 0 net17
rlabel metal1 2576 4114 2576 4114 0 net18
rlabel metal1 7590 7446 7590 7446 0 net2
rlabel metal1 8464 8942 8464 8942 0 net20
rlabel metal1 6394 7990 6394 7990 0 net21
rlabel metal1 1932 5678 1932 5678 0 net22
rlabel via1 3519 8942 3519 8942 0 net23
rlabel metal1 6440 4114 6440 4114 0 net24
rlabel metal1 1702 4590 1702 4590 0 net28
rlabel metal1 4600 4794 4600 4794 0 net3
rlabel metal1 1978 2618 1978 2618 0 net4
rlabel metal2 2070 9554 2070 9554 0 net5
rlabel metal2 3818 7548 3818 7548 0 net6
rlabel metal1 2484 7514 2484 7514 0 net7
rlabel metal1 5750 9622 5750 9622 0 net8
rlabel metal1 1840 9350 1840 9350 0 net9
rlabel metal1 8878 6766 8878 6766 0 reset
rlabel metal1 6854 9588 6854 9588 0 sel[0]
rlabel metal2 2070 2975 2070 2975 0 sel[1]
<< properties >>
string FIXED_BBOX 0 0 10212 12356
<< end >>
